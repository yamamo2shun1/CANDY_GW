-- candy_gw_qsys.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity candy_gw_qsys is
	port (
		adc_export                        : in    std_logic_vector(7 downto 0)  := (others => '0'); --                         adc.export
		altpll_locked_export              : out   std_logic;                                        --               altpll_locked.export
		clk_clk                           : in    std_logic                     := '0';             --                         clk.clk
		codec_clk_clk                     : out   std_logic;                                        --                   codec_clk.clk
		codec_reset_export                : out   std_logic;                                        --                 codec_reset.export
		grove1_in_port                    : in    std_logic_vector(1 downto 0)  := (others => '0'); --                      grove1.in_port
		grove1_out_port                   : out   std_logic_vector(1 downto 0);                     --                            .out_port
		i2s_lrclk_i_mst                   : in    std_logic                     := '0';             --                         i2s.lrclk_i_mst
		i2s_data_i_mst                    : in    std_logic                     := '0';             --                            .data_i_mst
		i2s_data_o_mst                    : out   std_logic;                                        --                            .data_o_mst
		i2s_lrclk_o_slv                   : out   std_logic;                                        --                            .lrclk_o_slv
		i2s_data_o_slv                    : out   std_logic;                                        --                            .data_o_slv
		i2s_bitclk_o_slv                  : out   std_logic;                                        --                            .bitclk_o_slv
		i2s_bclk_mst_clk                  : in    std_logic                     := '0';             --                i2s_bclk_mst.clk
		new_sdram_controller_0_wire_addr  : out   std_logic_vector(12 downto 0);                    -- new_sdram_controller_0_wire.addr
		new_sdram_controller_0_wire_ba    : out   std_logic_vector(1 downto 0);                     --                            .ba
		new_sdram_controller_0_wire_cas_n : out   std_logic;                                        --                            .cas_n
		new_sdram_controller_0_wire_cke   : out   std_logic;                                        --                            .cke
		new_sdram_controller_0_wire_cs_n  : out   std_logic;                                        --                            .cs_n
		new_sdram_controller_0_wire_dq    : inout std_logic_vector(15 downto 0) := (others => '0'); --                            .dq
		new_sdram_controller_0_wire_dqm   : out   std_logic_vector(1 downto 0);                     --                            .dqm
		new_sdram_controller_0_wire_ras_n : out   std_logic;                                        --                            .ras_n
		new_sdram_controller_0_wire_we_n  : out   std_logic;                                        --                            .we_n
		oe_export                         : out   std_logic;                                        --                          oe.export
		onbrd_led_pwm_out                 : out   std_logic_vector(3 downto 0);                     --                   onbrd_led.pwm_out
		pmod2_export                      : in    std_logic_vector(3 downto 0)  := (others => '0'); --                       pmod2.export
		qspi_dclk                         : out   std_logic;                                        --                        qspi.dclk
		qspi_ncs                          : out   std_logic;                                        --                            .ncs
		qspi_data                         : inout std_logic_vector(3 downto 0)  := (others => '0'); --                            .data
		reset_reset_n                     : in    std_logic                     := '0';             --                       reset.reset_n
		sdclk_clk_clk                     : out   std_logic;                                        --                   sdclk_clk.clk
		uart_rxd                          : in    std_logic                     := '0';             --                        uart.rxd
		uart_txd                          : out   std_logic;                                        --                            .txd
		uart_cts_n                        : in    std_logic                     := '0';             --                            .cts_n
		uart_rts_n                        : out   std_logic;                                        --                            .rts_n
		wb_ack_i                          : in    std_logic                     := '0';             --                          wb.ack_i
		wb_adr_o                          : out   std_logic_vector(31 downto 0);                    --                            .adr_o
		wb_clk_o                          : out   std_logic;                                        --                            .clk_o
		wb_cyc_o                          : out   std_logic;                                        --                            .cyc_o
		wb_dat_i                          : in    std_logic_vector(31 downto 0) := (others => '0'); --                            .dat_i
		wb_dat_o                          : out   std_logic_vector(31 downto 0);                    --                            .dat_o
		wb_err_i                          : in    std_logic                     := '0';             --                            .err_i
		wb_rst_o                          : out   std_logic;                                        --                            .rst_o
		wb_rty_i                          : in    std_logic                     := '0';             --                            .rty_i
		wb_sel_o                          : out   std_logic_vector(3 downto 0);                     --                            .sel_o
		wb_stb_o                          : out   std_logic;                                        --                            .stb_o
		wb_we_o                           : out   std_logic                                         --                            .we_o
	);
end entity candy_gw_qsys;

architecture rtl of candy_gw_qsys is
	component candy_gw_qsys_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component candy_gw_qsys_altpll_0;

	component AVALON_I2S is
		generic (
			DATA_WIDTH : integer := 32
		);
		port (
			csi_reset_n        : in  std_logic                     := 'X';             -- reset_n
			avs_s1_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avs_s1_write       : in  std_logic                     := 'X';             -- write
			avs_s1_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			LRCLK_I_MST        : in  std_logic                     := 'X';             -- lrclk_i_mst
			DATA_I_MST         : in  std_logic                     := 'X';             -- data_i_mst
			DATA_O_MST         : out std_logic;                                        -- data_o_mst
			LRCLK_O_SLV        : out std_logic;                                        -- lrclk_o_slv
			DATA_O_SLV         : out std_logic;                                        -- data_o_slv
			BITCLK_O_SLV       : out std_logic;                                        -- bitclk_o_slv
			av_mm2_address     : out std_logic_vector(2 downto 0);                     -- address
			av_mm2_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			av_mm2_read        : out std_logic;                                        -- read
			av_mm2_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_mm1_address     : out std_logic_vector(2 downto 0);                     -- address
			av_mm1_write       : out std_logic;                                        -- write
			av_mm1_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			av_mm1_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			bit_clk_mst        : in  std_logic                     := 'X'              -- clk
		);
	end component AVALON_I2S;

	component AVALON2PWM is
		generic (
			WIDTH           : integer := 3;
			PWM_COUNTER_MAX : integer := 60000
		);
		port (
			csi_clk          : in  std_logic                     := 'X';             -- clk
			csi_reset_n      : in  std_logic                     := 'X';             -- reset_n
			avs_s1_write     : in  std_logic                     := 'X';             -- write
			avs_s1_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s1_address   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avs_s1_read      : in  std_logic                     := 'X';             -- read
			avs_s1_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			PWM_OUT          : out std_logic_vector(3 downto 0)                      -- pwm_out
		);
	end component AVALON2PWM;

	component AVALON2WB is
		port (
			avs_s1_address       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avs_s1_chipselect    : in  std_logic                     := 'X';             -- chipselect
			avs_s1_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_s1_read          : in  std_logic                     := 'X';             -- read
			avs_s1_write         : in  std_logic                     := 'X';             -- write
			avs_s1_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s1_waitrequest   : out std_logic;                                        -- waitrequest
			avs_s1_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s1_readdatavalid : out std_logic;                                        -- readdatavalid
			ACK_I                : in  std_logic                     := 'X';             -- ack_i
			ADR_O                : out std_logic_vector(31 downto 0);                    -- adr_o
			CLK_O                : out std_logic;                                        -- clk_o
			CYC_O                : out std_logic;                                        -- cyc_o
			DAT_I                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dat_i
			DAT_O                : out std_logic_vector(31 downto 0);                    -- dat_o
			ERR_I                : in  std_logic                     := 'X';             -- err_i
			RST_O                : out std_logic;                                        -- rst_o
			RTY_I                : in  std_logic                     := 'X';             -- rty_i
			SEL_O                : out std_logic_vector(3 downto 0);                     -- sel_o
			STB_O                : out std_logic;                                        -- stb_o
			WE_O                 : out std_logic;                                        -- we_o
			csi_reset_n          : in  std_logic                     := 'X';             -- reset_n
			csi_clk              : in  std_logic                     := 'X'              -- clk
		);
	end component AVALON2WB;

	component candy_gw_qsys_dma_rx is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			system_reset_n     : in  std_logic                     := 'X';             -- reset_n
			dma_ctl_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			dma_ctl_chipselect : in  std_logic                     := 'X';             -- chipselect
			dma_ctl_readdata   : out std_logic_vector(24 downto 0);                    -- readdata
			dma_ctl_write_n    : in  std_logic                     := 'X';             -- write_n
			dma_ctl_writedata  : in  std_logic_vector(24 downto 0) := (others => 'X'); -- writedata
			dma_ctl_irq        : out std_logic;                                        -- irq
			read_address       : out std_logic_vector(4 downto 0);                     -- address
			read_chipselect    : out std_logic;                                        -- chipselect
			read_read_n        : out std_logic;                                        -- read_n
			read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			write_address      : out std_logic_vector(24 downto 0);                    -- address
			write_chipselect   : out std_logic;                                        -- chipselect
			write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			write_write_n      : out std_logic;                                        -- write_n
			write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			write_byteenable   : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component candy_gw_qsys_dma_rx;

	component candy_gw_qsys_dma_tx is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			system_reset_n     : in  std_logic                     := 'X';             -- reset_n
			dma_ctl_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			dma_ctl_chipselect : in  std_logic                     := 'X';             -- chipselect
			dma_ctl_readdata   : out std_logic_vector(24 downto 0);                    -- readdata
			dma_ctl_write_n    : in  std_logic                     := 'X';             -- write_n
			dma_ctl_writedata  : in  std_logic_vector(24 downto 0) := (others => 'X'); -- writedata
			dma_ctl_irq        : out std_logic;                                        -- irq
			read_address       : out std_logic_vector(24 downto 0);                    -- address
			read_chipselect    : out std_logic;                                        -- chipselect
			read_read_n        : out std_logic;                                        -- read_n
			read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			write_address      : out std_logic_vector(4 downto 0);                     -- address
			write_chipselect   : out std_logic;                                        -- chipselect
			write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			write_write_n      : out std_logic;                                        -- write_n
			write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			write_byteenable   : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component candy_gw_qsys_dma_tx;

	component candy_gw_qsys_fifo_rx is
		port (
			wrclock                        : in  std_logic                     := 'X';             -- clk
			reset_n                        : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write     : in  std_logic                     := 'X';             -- write
			avalonmm_read_slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read       : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read       : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write      : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			wrclk_control_slave_irq        : out std_logic                                         -- irq
		);
	end component candy_gw_qsys_fifo_rx;

	component candy_gw_qsys_fifo_tx is
		port (
			wrclock                        : in  std_logic                     := 'X';             -- clk
			reset_n                        : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write     : in  std_logic                     := 'X';             -- write
			avalonmm_read_slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read       : in  std_logic                     := 'X'              -- read
		);
	end component candy_gw_qsys_fifo_tx;

	component candy_gw_qsys_intel_generic_serial_flash_interface_top_0 is
		generic (
			DEVICE_FAMILY : string  := "";
			CHIP_SELS     : integer := 1
		);
		port (
			avl_csr_address       : in    std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			avl_csr_read          : in    std_logic                     := 'X';             -- read
			avl_csr_readdata      : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_csr_write         : in    std_logic                     := 'X';             -- write
			avl_csr_writedata     : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_csr_waitrequest   : out   std_logic;                                        -- waitrequest
			avl_csr_readdatavalid : out   std_logic;                                        -- readdatavalid
			avl_mem_write         : in    std_logic                     := 'X';             -- write
			avl_mem_burstcount    : in    std_logic_vector(6 downto 0)  := (others => 'X'); -- burstcount
			avl_mem_waitrequest   : out   std_logic;                                        -- waitrequest
			avl_mem_read          : in    std_logic                     := 'X';             -- read
			avl_mem_address       : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			avl_mem_writedata     : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_mem_readdata      : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_mem_readdatavalid : out   std_logic;                                        -- readdatavalid
			avl_mem_byteenable    : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk_clk               : in    std_logic                     := 'X';             -- clk
			reset_reset           : in    std_logic                     := 'X';             -- reset
			qspi_pins_dclk        : out   std_logic;                                        -- dclk
			qspi_pins_ncs         : out   std_logic;                                        -- ncs
			qspi_pins_data        : inout std_logic_vector(3 downto 0)  := (others => 'X')  -- data
		);
	end component candy_gw_qsys_intel_generic_serial_flash_interface_top_0;

	component candy_gw_qsys_jtaguart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component candy_gw_qsys_jtaguart_0;

	component candy_gw_qsys_new_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component candy_gw_qsys_new_sdram_controller_0;

	component candy_gw_qsys_nios2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			eic_port_valid                      : in  std_logic                     := 'X';             -- valid
			eic_port_data                       : in  std_logic_vector(44 downto 0) := (others => 'X'); -- data
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component candy_gw_qsys_nios2_0;

	component altera_onchip_flash is
		generic (
			INIT_FILENAME                       : string  := "";
			INIT_FILENAME_SIM                   : string  := "";
			DEVICE_FAMILY                       : string  := "Unknown";
			PART_NAME                           : string  := "Unknown";
			DEVICE_ID                           : string  := "Unknown";
			SECTOR1_START_ADDR                  : integer := 0;
			SECTOR1_END_ADDR                    : integer := 0;
			SECTOR2_START_ADDR                  : integer := 0;
			SECTOR2_END_ADDR                    : integer := 0;
			SECTOR3_START_ADDR                  : integer := 0;
			SECTOR3_END_ADDR                    : integer := 0;
			SECTOR4_START_ADDR                  : integer := 0;
			SECTOR4_END_ADDR                    : integer := 0;
			SECTOR5_START_ADDR                  : integer := 0;
			SECTOR5_END_ADDR                    : integer := 0;
			MIN_VALID_ADDR                      : integer := 0;
			MAX_VALID_ADDR                      : integer := 0;
			MIN_UFM_VALID_ADDR                  : integer := 0;
			MAX_UFM_VALID_ADDR                  : integer := 0;
			SECTOR1_MAP                         : integer := 0;
			SECTOR2_MAP                         : integer := 0;
			SECTOR3_MAP                         : integer := 0;
			SECTOR4_MAP                         : integer := 0;
			SECTOR5_MAP                         : integer := 0;
			ADDR_RANGE1_END_ADDR                : integer := 0;
			ADDR_RANGE2_END_ADDR                : integer := 0;
			ADDR_RANGE1_OFFSET                  : integer := 0;
			ADDR_RANGE2_OFFSET                  : integer := 0;
			ADDR_RANGE3_OFFSET                  : integer := 0;
			AVMM_DATA_ADDR_WIDTH                : integer := 19;
			AVMM_DATA_DATA_WIDTH                : integer := 32;
			AVMM_DATA_BURSTCOUNT_WIDTH          : integer := 4;
			SECTOR_READ_PROTECTION_MODE         : integer := 31;
			FLASH_SEQ_READ_DATA_COUNT           : integer := 2;
			FLASH_ADDR_ALIGNMENT_BITS           : integer := 1;
			FLASH_READ_CYCLE_MAX_INDEX          : integer := 4;
			FLASH_RESET_CYCLE_MAX_INDEX         : integer := 29;
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  : integer := 112;
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX : integer := 40603248;
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX : integer := 35382;
			PARALLEL_MODE                       : boolean := true;
			READ_AND_WRITE_MODE                 : boolean := true;
			WRAPPING_BURST_MODE                 : boolean := false;
			IS_DUAL_BOOT                        : string  := "False";
			IS_ERAM_SKIP                        : string  := "False";
			IS_COMPRESSED_IMAGE                 : string  := "False"
		);
		port (
			clock                   : in  std_logic                     := 'X';             -- clk
			reset_n                 : in  std_logic                     := 'X';             -- reset_n
			avmm_data_addr          : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			avmm_data_read          : in  std_logic                     := 'X';             -- read
			avmm_data_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_data_write         : in  std_logic                     := 'X';             -- write
			avmm_data_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avmm_data_waitrequest   : out std_logic;                                        -- waitrequest
			avmm_data_readdatavalid : out std_logic;                                        -- readdatavalid
			avmm_data_burstcount    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			avmm_csr_addr           : in  std_logic                     := 'X';             -- address
			avmm_csr_read           : in  std_logic                     := 'X';             -- read
			avmm_csr_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_csr_write          : in  std_logic                     := 'X';             -- write
			avmm_csr_readdata       : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component altera_onchip_flash;

	component candy_gw_qsys_pio_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component candy_gw_qsys_pio_1;

	component candy_gw_qsys_pio_3 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component candy_gw_qsys_pio_3;

	component candy_gw_qsys_pio_4 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component candy_gw_qsys_pio_4;

	component candy_gw_qsys_pio_6 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component candy_gw_qsys_pio_6;

	component candy_gw_qsys_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component candy_gw_qsys_sys_clk_timer;

	component candy_gw_qsys_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component candy_gw_qsys_sysid;

	component candy_gw_qsys_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component candy_gw_qsys_timer_0;

	component candy_gw_qsys_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			cts_n         : in  std_logic                     := 'X';             -- export
			rts_n         : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component candy_gw_qsys_uart_0;

	component candy_gw_qsys_vic_0 is
		port (
			clk_clk                        : in  std_logic                     := 'X';             -- clk
			reset_reset                    : in  std_logic                     := 'X';             -- reset
			irq_input_irq                  : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- irq
			csr_access_read                : in  std_logic                     := 'X';             -- read
			csr_access_write               : in  std_logic                     := 'X';             -- write
			csr_access_address             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			csr_access_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_access_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			interrupt_controller_out_valid : out std_logic;                                        -- valid
			interrupt_controller_out_data  : out std_logic_vector(44 downto 0)                     -- data
		);
	end component candy_gw_qsys_vic_0;

	component candy_gw_qsys_mm_interconnect_0 is
		port (
			altpll_0_c1_clk                                : in  std_logic                     := 'X';             -- clk
			clock_bridge_0_out_clk_clk                     : in  std_logic                     := 'X';             -- clk
			avalon_i2s_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			fifo_rx_reset_in_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			avalon_i2s_0_av_mm1_address                    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avalon_i2s_0_av_mm1_waitrequest                : out std_logic;                                        -- waitrequest
			avalon_i2s_0_av_mm1_write                      : in  std_logic                     := 'X';             -- write
			avalon_i2s_0_av_mm1_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			fifo_rx_in_write                               : out std_logic;                                        -- write
			fifo_rx_in_writedata                           : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component candy_gw_qsys_mm_interconnect_0;

	component candy_gw_qsys_mm_interconnect_1 is
		port (
			altpll_0_c1_clk                                : in  std_logic                     := 'X';             -- clk
			clock_bridge_0_out_clk_clk                     : in  std_logic                     := 'X';             -- clk
			avalon_i2s_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			fifo_tx_reset_in_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			avalon_i2s_0_av_mm2_address                    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avalon_i2s_0_av_mm2_waitrequest                : out std_logic;                                        -- waitrequest
			avalon_i2s_0_av_mm2_read                       : in  std_logic                     := 'X';             -- read
			avalon_i2s_0_av_mm2_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			fifo_tx_out_read                               : out std_logic;                                        -- read
			fifo_tx_out_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component candy_gw_qsys_mm_interconnect_1;

	component candy_gw_qsys_mm_interconnect_2 is
		port (
			altpll_0_c1_clk                                                              : in  std_logic                     := 'X';             -- clk
			clk_0_clk_clk                                                                : in  std_logic                     := 'X';             -- clk
			clock_bridge_0_out_clk_clk                                                   : in  std_logic                     := 'X';             -- clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset                   : in  std_logic                     := 'X';             -- reset
			avalon_i2s_0_reset_reset_bridge_in_reset_reset                               : in  std_logic                     := 'X';             -- reset
			intel_generic_serial_flash_interface_top_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_0_reset_reset_bridge_in_reset_reset                                    : in  std_logic                     := 'X';             -- reset
			dma_rx_write_master_address                                                  : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			dma_rx_write_master_waitrequest                                              : out std_logic;                                        -- waitrequest
			dma_rx_write_master_byteenable                                               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			dma_rx_write_master_chipselect                                               : in  std_logic                     := 'X';             -- chipselect
			dma_rx_write_master_write                                                    : in  std_logic                     := 'X';             -- write
			dma_rx_write_master_writedata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dma_tx_read_master_address                                                   : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			dma_tx_read_master_waitrequest                                               : out std_logic;                                        -- waitrequest
			dma_tx_read_master_chipselect                                                : in  std_logic                     := 'X';             -- chipselect
			dma_tx_read_master_read                                                      : in  std_logic                     := 'X';             -- read
			dma_tx_read_master_readdata                                                  : out std_logic_vector(31 downto 0);                    -- readdata
			dma_tx_read_master_readdatavalid                                             : out std_logic;                                        -- readdatavalid
			nios2_0_data_master_address                                                  : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_0_data_master_waitrequest                                              : out std_logic;                                        -- waitrequest
			nios2_0_data_master_byteenable                                               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_0_data_master_read                                                     : in  std_logic                     := 'X';             -- read
			nios2_0_data_master_readdata                                                 : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_0_data_master_readdatavalid                                            : out std_logic;                                        -- readdatavalid
			nios2_0_data_master_write                                                    : in  std_logic                     := 'X';             -- write
			nios2_0_data_master_writedata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_0_data_master_debugaccess                                              : in  std_logic                     := 'X';             -- debugaccess
			nios2_0_instruction_master_address                                           : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_0_instruction_master_waitrequest                                       : out std_logic;                                        -- waitrequest
			nios2_0_instruction_master_read                                              : in  std_logic                     := 'X';             -- read
			nios2_0_instruction_master_readdata                                          : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_0_instruction_master_readdatavalid                                     : out std_logic;                                        -- readdatavalid
			altpll_0_pll_slave_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                                     : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                                      : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			avalon_i2s_0_s1_address                                                      : out std_logic_vector(1 downto 0);                     -- address
			avalon_i2s_0_s1_write                                                        : out std_logic;                                        -- write
			avalon_i2s_0_s1_writedata                                                    : out std_logic_vector(31 downto 0);                    -- writedata
			avalon_pwm_0_s1_address                                                      : out std_logic_vector(2 downto 0);                     -- address
			avalon_pwm_0_s1_write                                                        : out std_logic;                                        -- write
			avalon_pwm_0_s1_read                                                         : out std_logic;                                        -- read
			avalon_pwm_0_s1_readdata                                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avalon_pwm_0_s1_writedata                                                    : out std_logic_vector(31 downto 0);                    -- writedata
			avalon_wb_s1_address                                                         : out std_logic_vector(7 downto 0);                     -- address
			avalon_wb_s1_write                                                           : out std_logic;                                        -- write
			avalon_wb_s1_read                                                            : out std_logic;                                        -- read
			avalon_wb_s1_readdata                                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avalon_wb_s1_writedata                                                       : out std_logic_vector(31 downto 0);                    -- writedata
			avalon_wb_s1_byteenable                                                      : out std_logic_vector(3 downto 0);                     -- byteenable
			avalon_wb_s1_readdatavalid                                                   : in  std_logic                     := 'X';             -- readdatavalid
			avalon_wb_s1_waitrequest                                                     : in  std_logic                     := 'X';             -- waitrequest
			avalon_wb_s1_chipselect                                                      : out std_logic;                                        -- chipselect
			dma_rx_control_port_slave_address                                            : out std_logic_vector(2 downto 0);                     -- address
			dma_rx_control_port_slave_write                                              : out std_logic;                                        -- write
			dma_rx_control_port_slave_readdata                                           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- readdata
			dma_rx_control_port_slave_writedata                                          : out std_logic_vector(24 downto 0);                    -- writedata
			dma_rx_control_port_slave_chipselect                                         : out std_logic;                                        -- chipselect
			dma_tx_control_port_slave_address                                            : out std_logic_vector(2 downto 0);                     -- address
			dma_tx_control_port_slave_write                                              : out std_logic;                                        -- write
			dma_tx_control_port_slave_readdata                                           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- readdata
			dma_tx_control_port_slave_writedata                                          : out std_logic_vector(24 downto 0);                    -- writedata
			dma_tx_control_port_slave_chipselect                                         : out std_logic;                                        -- chipselect
			fifo_rx_in_csr_address                                                       : out std_logic_vector(2 downto 0);                     -- address
			fifo_rx_in_csr_write                                                         : out std_logic;                                        -- write
			fifo_rx_in_csr_read                                                          : out std_logic;                                        -- read
			fifo_rx_in_csr_readdata                                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_rx_in_csr_writedata                                                     : out std_logic_vector(31 downto 0);                    -- writedata
			intel_generic_serial_flash_interface_top_0_avl_csr_address                   : out std_logic_vector(5 downto 0);                     -- address
			intel_generic_serial_flash_interface_top_0_avl_csr_write                     : out std_logic;                                        -- write
			intel_generic_serial_flash_interface_top_0_avl_csr_read                      : out std_logic;                                        -- read
			intel_generic_serial_flash_interface_top_0_avl_csr_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			intel_generic_serial_flash_interface_top_0_avl_csr_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid             : in  std_logic                     := 'X';             -- readdatavalid
			intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			intel_generic_serial_flash_interface_top_0_avl_mem_address                   : out std_logic_vector(21 downto 0);                    -- address
			intel_generic_serial_flash_interface_top_0_avl_mem_write                     : out std_logic;                                        -- write
			intel_generic_serial_flash_interface_top_0_avl_mem_read                      : out std_logic;                                        -- read
			intel_generic_serial_flash_interface_top_0_avl_mem_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			intel_generic_serial_flash_interface_top_0_avl_mem_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			intel_generic_serial_flash_interface_top_0_avl_mem_burstcount                : out std_logic_vector(6 downto 0);                     -- burstcount
			intel_generic_serial_flash_interface_top_0_avl_mem_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid             : in  std_logic                     := 'X';             -- readdatavalid
			intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtaguart_0_avalon_jtag_slave_address                                         : out std_logic_vector(0 downto 0);                     -- address
			jtaguart_0_avalon_jtag_slave_write                                           : out std_logic;                                        -- write
			jtaguart_0_avalon_jtag_slave_read                                            : out std_logic;                                        -- read
			jtaguart_0_avalon_jtag_slave_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtaguart_0_avalon_jtag_slave_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			jtaguart_0_avalon_jtag_slave_waitrequest                                     : in  std_logic                     := 'X';             -- waitrequest
			jtaguart_0_avalon_jtag_slave_chipselect                                      : out std_logic;                                        -- chipselect
			new_sdram_controller_0_s1_address                                            : out std_logic_vector(23 downto 0);                    -- address
			new_sdram_controller_0_s1_write                                              : out std_logic;                                        -- write
			new_sdram_controller_0_s1_read                                               : out std_logic;                                        -- read
			new_sdram_controller_0_s1_readdata                                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			new_sdram_controller_0_s1_writedata                                          : out std_logic_vector(15 downto 0);                    -- writedata
			new_sdram_controller_0_s1_byteenable                                         : out std_logic_vector(1 downto 0);                     -- byteenable
			new_sdram_controller_0_s1_readdatavalid                                      : in  std_logic                     := 'X';             -- readdatavalid
			new_sdram_controller_0_s1_waitrequest                                        : in  std_logic                     := 'X';             -- waitrequest
			new_sdram_controller_0_s1_chipselect                                         : out std_logic;                                        -- chipselect
			nios2_0_debug_mem_slave_address                                              : out std_logic_vector(8 downto 0);                     -- address
			nios2_0_debug_mem_slave_write                                                : out std_logic;                                        -- write
			nios2_0_debug_mem_slave_read                                                 : out std_logic;                                        -- read
			nios2_0_debug_mem_slave_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_0_debug_mem_slave_writedata                                            : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_0_debug_mem_slave_byteenable                                           : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_0_debug_mem_slave_waitrequest                                          : in  std_logic                     := 'X';             -- waitrequest
			nios2_0_debug_mem_slave_debugaccess                                          : out std_logic;                                        -- debugaccess
			onchip_flash_0_csr_address                                                   : out std_logic_vector(0 downto 0);                     -- address
			onchip_flash_0_csr_write                                                     : out std_logic;                                        -- write
			onchip_flash_0_csr_read                                                      : out std_logic;                                        -- read
			onchip_flash_0_csr_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_0_csr_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_0_data_address                                                  : out std_logic_vector(17 downto 0);                    -- address
			onchip_flash_0_data_write                                                    : out std_logic;                                        -- write
			onchip_flash_0_data_read                                                     : out std_logic;                                        -- read
			onchip_flash_0_data_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_0_data_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_0_data_burstcount                                               : out std_logic_vector(3 downto 0);                     -- burstcount
			onchip_flash_0_data_readdatavalid                                            : in  std_logic                     := 'X';             -- readdatavalid
			onchip_flash_0_data_waitrequest                                              : in  std_logic                     := 'X';             -- waitrequest
			pio_1_s1_address                                                             : out std_logic_vector(1 downto 0);                     -- address
			pio_1_s1_write                                                               : out std_logic;                                        -- write
			pio_1_s1_readdata                                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_1_s1_writedata                                                           : out std_logic_vector(31 downto 0);                    -- writedata
			pio_1_s1_chipselect                                                          : out std_logic;                                        -- chipselect
			pio_3_s1_address                                                             : out std_logic_vector(1 downto 0);                     -- address
			pio_3_s1_readdata                                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_4_s1_address                                                             : out std_logic_vector(1 downto 0);                     -- address
			pio_4_s1_write                                                               : out std_logic;                                        -- write
			pio_4_s1_readdata                                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_4_s1_writedata                                                           : out std_logic_vector(31 downto 0);                    -- writedata
			pio_4_s1_chipselect                                                          : out std_logic;                                        -- chipselect
			pio_5_s1_address                                                             : out std_logic_vector(1 downto 0);                     -- address
			pio_5_s1_write                                                               : out std_logic;                                        -- write
			pio_5_s1_readdata                                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_5_s1_writedata                                                           : out std_logic_vector(31 downto 0);                    -- writedata
			pio_5_s1_chipselect                                                          : out std_logic;                                        -- chipselect
			pio_6_s1_address                                                             : out std_logic_vector(1 downto 0);                     -- address
			pio_6_s1_readdata                                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_address                                                     : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                                                       : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata                                                    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata                                                   : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect                                                  : out std_logic;                                        -- chipselect
			sysid_control_slave_address                                                  : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                                           : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                                             : out std_logic;                                        -- write
			timer_0_s1_readdata                                                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                                         : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                                        : out std_logic;                                        -- chipselect
			uart_0_s1_address                                                            : out std_logic_vector(2 downto 0);                     -- address
			uart_0_s1_write                                                              : out std_logic;                                        -- write
			uart_0_s1_read                                                               : out std_logic;                                        -- read
			uart_0_s1_readdata                                                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_0_s1_writedata                                                          : out std_logic_vector(15 downto 0);                    -- writedata
			uart_0_s1_begintransfer                                                      : out std_logic;                                        -- begintransfer
			uart_0_s1_chipselect                                                         : out std_logic;                                        -- chipselect
			vic_0_csr_access_address                                                     : out std_logic_vector(7 downto 0);                     -- address
			vic_0_csr_access_write                                                       : out std_logic;                                        -- write
			vic_0_csr_access_read                                                        : out std_logic;                                        -- read
			vic_0_csr_access_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vic_0_csr_access_writedata                                                   : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component candy_gw_qsys_mm_interconnect_2;

	component candy_gw_qsys_mm_interconnect_3 is
		port (
			altpll_0_c1_clk                          : in  std_logic                     := 'X';             -- clk
			dma_rx_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			dma_rx_read_master_address               : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			dma_rx_read_master_waitrequest           : out std_logic;                                        -- waitrequest
			dma_rx_read_master_chipselect            : in  std_logic                     := 'X';             -- chipselect
			dma_rx_read_master_read                  : in  std_logic                     := 'X';             -- read
			dma_rx_read_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			dma_rx_read_master_readdatavalid         : out std_logic;                                        -- readdatavalid
			fifo_rx_out_read                         : out std_logic;                                        -- read
			fifo_rx_out_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component candy_gw_qsys_mm_interconnect_3;

	component candy_gw_qsys_mm_interconnect_4 is
		port (
			altpll_0_c1_clk                          : in  std_logic                     := 'X';             -- clk
			dma_tx_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			dma_tx_write_master_address              : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			dma_tx_write_master_waitrequest          : out std_logic;                                        -- waitrequest
			dma_tx_write_master_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			dma_tx_write_master_chipselect           : in  std_logic                     := 'X';             -- chipselect
			dma_tx_write_master_write                : in  std_logic                     := 'X';             -- write
			dma_tx_write_master_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			fifo_tx_in_write                         : out std_logic;                                        -- write
			fifo_tx_in_writedata                     : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component candy_gw_qsys_mm_interconnect_4;

	component candy_gw_qsys_irq_mapper is
		port (
			clk           : in  std_logic                    := 'X'; -- clk
			reset         : in  std_logic                    := 'X'; -- reset
			receiver0_irq : in  std_logic                    := 'X'; -- irq
			receiver1_irq : in  std_logic                    := 'X'; -- irq
			receiver2_irq : in  std_logic                    := 'X'; -- irq
			receiver3_irq : in  std_logic                    := 'X'; -- irq
			receiver4_irq : in  std_logic                    := 'X'; -- irq
			receiver5_irq : in  std_logic                    := 'X'; -- irq
			receiver6_irq : in  std_logic                    := 'X'; -- irq
			sender_irq    : out std_logic_vector(6 downto 0)         -- irq
		);
	end component candy_gw_qsys_irq_mapper;

	component candy_gw_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component candy_gw_qsys_rst_controller;

	component candy_gw_qsys_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component candy_gw_qsys_rst_controller_002;

	signal vic_0_interrupt_controller_out_valid                                               : std_logic;                     -- vic_0:interrupt_controller_out_valid -> nios2_0:eic_port_valid
	signal vic_0_interrupt_controller_out_data                                                : std_logic_vector(44 downto 0); -- vic_0:interrupt_controller_out_data -> nios2_0:eic_port_data
	signal altpll_0_c1_clk                                                                    : std_logic;                     -- altpll_0:c1 -> [avalon_pwm_0:csi_clk, avalon_wb:csi_clk, dma_rx:clk, dma_tx:clk, fifo_rx:wrclock, fifo_tx:wrclock, intel_generic_serial_flash_interface_top_0:clk_clk, irq_mapper:clk, jtaguart_0:clk, mm_interconnect_0:altpll_0_c1_clk, mm_interconnect_1:altpll_0_c1_clk, mm_interconnect_2:altpll_0_c1_clk, mm_interconnect_3:altpll_0_c1_clk, mm_interconnect_4:altpll_0_c1_clk, new_sdram_controller_0:clk, nios2_0:clk, onchip_flash_0:clock, pio_1:clk, pio_3:clk, pio_4:clk, pio_5:clk, pio_6:clk, rst_controller_002:clk, sys_clk_timer:clk, sysid:clock, timer_0:clk, uart_0:clk, vic_0:clk_clk]
	signal avalon_i2s_0_av_mm1_waitrequest                                                    : std_logic;                     -- mm_interconnect_0:avalon_i2s_0_av_mm1_waitrequest -> avalon_i2s_0:av_mm1_waitrequest
	signal avalon_i2s_0_av_mm1_address                                                        : std_logic_vector(2 downto 0);  -- avalon_i2s_0:av_mm1_address -> mm_interconnect_0:avalon_i2s_0_av_mm1_address
	signal avalon_i2s_0_av_mm1_write                                                          : std_logic;                     -- avalon_i2s_0:av_mm1_write -> mm_interconnect_0:avalon_i2s_0_av_mm1_write
	signal avalon_i2s_0_av_mm1_writedata                                                      : std_logic_vector(31 downto 0); -- avalon_i2s_0:av_mm1_writedata -> mm_interconnect_0:avalon_i2s_0_av_mm1_writedata
	signal mm_interconnect_0_fifo_rx_in_write                                                 : std_logic;                     -- mm_interconnect_0:fifo_rx_in_write -> fifo_rx:avalonmm_write_slave_write
	signal mm_interconnect_0_fifo_rx_in_writedata                                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:fifo_rx_in_writedata -> fifo_rx:avalonmm_write_slave_writedata
	signal avalon_i2s_0_av_mm2_waitrequest                                                    : std_logic;                     -- mm_interconnect_1:avalon_i2s_0_av_mm2_waitrequest -> avalon_i2s_0:av_mm2_waitrequest
	signal avalon_i2s_0_av_mm2_readdata                                                       : std_logic_vector(31 downto 0); -- mm_interconnect_1:avalon_i2s_0_av_mm2_readdata -> avalon_i2s_0:av_mm2_readdata
	signal avalon_i2s_0_av_mm2_address                                                        : std_logic_vector(2 downto 0);  -- avalon_i2s_0:av_mm2_address -> mm_interconnect_1:avalon_i2s_0_av_mm2_address
	signal avalon_i2s_0_av_mm2_read                                                           : std_logic;                     -- avalon_i2s_0:av_mm2_read -> mm_interconnect_1:avalon_i2s_0_av_mm2_read
	signal mm_interconnect_1_fifo_tx_out_readdata                                             : std_logic_vector(31 downto 0); -- fifo_tx:avalonmm_read_slave_readdata -> mm_interconnect_1:fifo_tx_out_readdata
	signal mm_interconnect_1_fifo_tx_out_read                                                 : std_logic;                     -- mm_interconnect_1:fifo_tx_out_read -> fifo_tx:avalonmm_read_slave_read
	signal nios2_0_data_master_readdata                                                       : std_logic_vector(31 downto 0); -- mm_interconnect_2:nios2_0_data_master_readdata -> nios2_0:d_readdata
	signal nios2_0_data_master_waitrequest                                                    : std_logic;                     -- mm_interconnect_2:nios2_0_data_master_waitrequest -> nios2_0:d_waitrequest
	signal nios2_0_data_master_debugaccess                                                    : std_logic;                     -- nios2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_2:nios2_0_data_master_debugaccess
	signal nios2_0_data_master_address                                                        : std_logic_vector(26 downto 0); -- nios2_0:d_address -> mm_interconnect_2:nios2_0_data_master_address
	signal nios2_0_data_master_byteenable                                                     : std_logic_vector(3 downto 0);  -- nios2_0:d_byteenable -> mm_interconnect_2:nios2_0_data_master_byteenable
	signal nios2_0_data_master_read                                                           : std_logic;                     -- nios2_0:d_read -> mm_interconnect_2:nios2_0_data_master_read
	signal nios2_0_data_master_readdatavalid                                                  : std_logic;                     -- mm_interconnect_2:nios2_0_data_master_readdatavalid -> nios2_0:d_readdatavalid
	signal nios2_0_data_master_write                                                          : std_logic;                     -- nios2_0:d_write -> mm_interconnect_2:nios2_0_data_master_write
	signal nios2_0_data_master_writedata                                                      : std_logic_vector(31 downto 0); -- nios2_0:d_writedata -> mm_interconnect_2:nios2_0_data_master_writedata
	signal nios2_0_instruction_master_readdata                                                : std_logic_vector(31 downto 0); -- mm_interconnect_2:nios2_0_instruction_master_readdata -> nios2_0:i_readdata
	signal nios2_0_instruction_master_waitrequest                                             : std_logic;                     -- mm_interconnect_2:nios2_0_instruction_master_waitrequest -> nios2_0:i_waitrequest
	signal nios2_0_instruction_master_address                                                 : std_logic_vector(26 downto 0); -- nios2_0:i_address -> mm_interconnect_2:nios2_0_instruction_master_address
	signal nios2_0_instruction_master_read                                                    : std_logic;                     -- nios2_0:i_read -> mm_interconnect_2:nios2_0_instruction_master_read
	signal nios2_0_instruction_master_readdatavalid                                           : std_logic;                     -- mm_interconnect_2:nios2_0_instruction_master_readdatavalid -> nios2_0:i_readdatavalid
	signal dma_tx_read_master_chipselect                                                      : std_logic;                     -- dma_tx:read_chipselect -> mm_interconnect_2:dma_tx_read_master_chipselect
	signal dma_tx_read_master_readdata                                                        : std_logic_vector(31 downto 0); -- mm_interconnect_2:dma_tx_read_master_readdata -> dma_tx:read_readdata
	signal dma_tx_read_master_waitrequest                                                     : std_logic;                     -- mm_interconnect_2:dma_tx_read_master_waitrequest -> dma_tx:read_waitrequest
	signal dma_tx_read_master_address                                                         : std_logic_vector(24 downto 0); -- dma_tx:read_address -> mm_interconnect_2:dma_tx_read_master_address
	signal dma_tx_read_master_read                                                            : std_logic;                     -- dma_tx:read_read_n -> dma_tx_read_master_read:in
	signal dma_tx_read_master_readdatavalid                                                   : std_logic;                     -- mm_interconnect_2:dma_tx_read_master_readdatavalid -> dma_tx:read_readdatavalid
	signal dma_rx_write_master_chipselect                                                     : std_logic;                     -- dma_rx:write_chipselect -> mm_interconnect_2:dma_rx_write_master_chipselect
	signal dma_rx_write_master_waitrequest                                                    : std_logic;                     -- mm_interconnect_2:dma_rx_write_master_waitrequest -> dma_rx:write_waitrequest
	signal dma_rx_write_master_address                                                        : std_logic_vector(24 downto 0); -- dma_rx:write_address -> mm_interconnect_2:dma_rx_write_master_address
	signal dma_rx_write_master_byteenable                                                     : std_logic_vector(3 downto 0);  -- dma_rx:write_byteenable -> mm_interconnect_2:dma_rx_write_master_byteenable
	signal dma_rx_write_master_write                                                          : std_logic;                     -- dma_rx:write_write_n -> dma_rx_write_master_write:in
	signal dma_rx_write_master_writedata                                                      : std_logic_vector(31 downto 0); -- dma_rx:write_writedata -> mm_interconnect_2:dma_rx_write_master_writedata
	signal mm_interconnect_2_jtaguart_0_avalon_jtag_slave_chipselect                          : std_logic;                     -- mm_interconnect_2:jtaguart_0_avalon_jtag_slave_chipselect -> jtaguart_0:av_chipselect
	signal mm_interconnect_2_jtaguart_0_avalon_jtag_slave_readdata                            : std_logic_vector(31 downto 0); -- jtaguart_0:av_readdata -> mm_interconnect_2:jtaguart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_2_jtaguart_0_avalon_jtag_slave_waitrequest                         : std_logic;                     -- jtaguart_0:av_waitrequest -> mm_interconnect_2:jtaguart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_2_jtaguart_0_avalon_jtag_slave_address                             : std_logic_vector(0 downto 0);  -- mm_interconnect_2:jtaguart_0_avalon_jtag_slave_address -> jtaguart_0:av_address
	signal mm_interconnect_2_jtaguart_0_avalon_jtag_slave_read                                : std_logic;                     -- mm_interconnect_2:jtaguart_0_avalon_jtag_slave_read -> mm_interconnect_2_jtaguart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_2_jtaguart_0_avalon_jtag_slave_write                               : std_logic;                     -- mm_interconnect_2:jtaguart_0_avalon_jtag_slave_write -> mm_interconnect_2_jtaguart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_2_jtaguart_0_avalon_jtag_slave_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_2:jtaguart_0_avalon_jtag_slave_writedata -> jtaguart_0:av_writedata
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_readdata      : std_logic_vector(31 downto 0); -- intel_generic_serial_flash_interface_top_0:avl_csr_readdata -> mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_csr_readdata
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest   : std_logic;                     -- intel_generic_serial_flash_interface_top_0:avl_csr_waitrequest -> mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_address       : std_logic_vector(5 downto 0);  -- mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_csr_address -> intel_generic_serial_flash_interface_top_0:avl_csr_address
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_read          : std_logic;                     -- mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_csr_read -> intel_generic_serial_flash_interface_top_0:avl_csr_read
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid : std_logic;                     -- intel_generic_serial_flash_interface_top_0:avl_csr_readdatavalid -> mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_write         : std_logic;                     -- mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_csr_write -> intel_generic_serial_flash_interface_top_0:avl_csr_write
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_csr_writedata -> intel_generic_serial_flash_interface_top_0:avl_csr_writedata
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_readdata      : std_logic_vector(31 downto 0); -- intel_generic_serial_flash_interface_top_0:avl_mem_readdata -> mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_mem_readdata
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest   : std_logic;                     -- intel_generic_serial_flash_interface_top_0:avl_mem_waitrequest -> mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_address       : std_logic_vector(21 downto 0); -- mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_mem_address -> intel_generic_serial_flash_interface_top_0:avl_mem_address
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_read          : std_logic;                     -- mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_mem_read -> intel_generic_serial_flash_interface_top_0:avl_mem_read
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_mem_byteenable -> intel_generic_serial_flash_interface_top_0:avl_mem_byteenable
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid : std_logic;                     -- intel_generic_serial_flash_interface_top_0:avl_mem_readdatavalid -> mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_write         : std_logic;                     -- mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_mem_write -> intel_generic_serial_flash_interface_top_0:avl_mem_write
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_mem_writedata -> intel_generic_serial_flash_interface_top_0:avl_mem_writedata
	signal mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_burstcount    : std_logic_vector(6 downto 0);  -- mm_interconnect_2:intel_generic_serial_flash_interface_top_0_avl_mem_burstcount -> intel_generic_serial_flash_interface_top_0:avl_mem_burstcount
	signal mm_interconnect_2_dma_rx_control_port_slave_chipselect                             : std_logic;                     -- mm_interconnect_2:dma_rx_control_port_slave_chipselect -> dma_rx:dma_ctl_chipselect
	signal mm_interconnect_2_dma_rx_control_port_slave_readdata                               : std_logic_vector(24 downto 0); -- dma_rx:dma_ctl_readdata -> mm_interconnect_2:dma_rx_control_port_slave_readdata
	signal mm_interconnect_2_dma_rx_control_port_slave_address                                : std_logic_vector(2 downto 0);  -- mm_interconnect_2:dma_rx_control_port_slave_address -> dma_rx:dma_ctl_address
	signal mm_interconnect_2_dma_rx_control_port_slave_write                                  : std_logic;                     -- mm_interconnect_2:dma_rx_control_port_slave_write -> mm_interconnect_2_dma_rx_control_port_slave_write:in
	signal mm_interconnect_2_dma_rx_control_port_slave_writedata                              : std_logic_vector(24 downto 0); -- mm_interconnect_2:dma_rx_control_port_slave_writedata -> dma_rx:dma_ctl_writedata
	signal mm_interconnect_2_dma_tx_control_port_slave_chipselect                             : std_logic;                     -- mm_interconnect_2:dma_tx_control_port_slave_chipselect -> dma_tx:dma_ctl_chipselect
	signal mm_interconnect_2_dma_tx_control_port_slave_readdata                               : std_logic_vector(24 downto 0); -- dma_tx:dma_ctl_readdata -> mm_interconnect_2:dma_tx_control_port_slave_readdata
	signal mm_interconnect_2_dma_tx_control_port_slave_address                                : std_logic_vector(2 downto 0);  -- mm_interconnect_2:dma_tx_control_port_slave_address -> dma_tx:dma_ctl_address
	signal mm_interconnect_2_dma_tx_control_port_slave_write                                  : std_logic;                     -- mm_interconnect_2:dma_tx_control_port_slave_write -> mm_interconnect_2_dma_tx_control_port_slave_write:in
	signal mm_interconnect_2_dma_tx_control_port_slave_writedata                              : std_logic_vector(24 downto 0); -- mm_interconnect_2:dma_tx_control_port_slave_writedata -> dma_tx:dma_ctl_writedata
	signal mm_interconnect_2_sysid_control_slave_readdata                                     : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_2:sysid_control_slave_readdata
	signal mm_interconnect_2_sysid_control_slave_address                                      : std_logic_vector(0 downto 0);  -- mm_interconnect_2:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_2_onchip_flash_0_csr_readdata                                      : std_logic_vector(31 downto 0); -- onchip_flash_0:avmm_csr_readdata -> mm_interconnect_2:onchip_flash_0_csr_readdata
	signal mm_interconnect_2_onchip_flash_0_csr_address                                       : std_logic_vector(0 downto 0);  -- mm_interconnect_2:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	signal mm_interconnect_2_onchip_flash_0_csr_read                                          : std_logic;                     -- mm_interconnect_2:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	signal mm_interconnect_2_onchip_flash_0_csr_write                                         : std_logic;                     -- mm_interconnect_2:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	signal mm_interconnect_2_onchip_flash_0_csr_writedata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_2:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	signal mm_interconnect_2_vic_0_csr_access_readdata                                        : std_logic_vector(31 downto 0); -- vic_0:csr_access_readdata -> mm_interconnect_2:vic_0_csr_access_readdata
	signal mm_interconnect_2_vic_0_csr_access_address                                         : std_logic_vector(7 downto 0);  -- mm_interconnect_2:vic_0_csr_access_address -> vic_0:csr_access_address
	signal mm_interconnect_2_vic_0_csr_access_read                                            : std_logic;                     -- mm_interconnect_2:vic_0_csr_access_read -> vic_0:csr_access_read
	signal mm_interconnect_2_vic_0_csr_access_write                                           : std_logic;                     -- mm_interconnect_2:vic_0_csr_access_write -> vic_0:csr_access_write
	signal mm_interconnect_2_vic_0_csr_access_writedata                                       : std_logic_vector(31 downto 0); -- mm_interconnect_2:vic_0_csr_access_writedata -> vic_0:csr_access_writedata
	signal mm_interconnect_2_onchip_flash_0_data_readdata                                     : std_logic_vector(31 downto 0); -- onchip_flash_0:avmm_data_readdata -> mm_interconnect_2:onchip_flash_0_data_readdata
	signal mm_interconnect_2_onchip_flash_0_data_waitrequest                                  : std_logic;                     -- onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_2:onchip_flash_0_data_waitrequest
	signal mm_interconnect_2_onchip_flash_0_data_address                                      : std_logic_vector(17 downto 0); -- mm_interconnect_2:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	signal mm_interconnect_2_onchip_flash_0_data_read                                         : std_logic;                     -- mm_interconnect_2:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	signal mm_interconnect_2_onchip_flash_0_data_readdatavalid                                : std_logic;                     -- onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_2:onchip_flash_0_data_readdatavalid
	signal mm_interconnect_2_onchip_flash_0_data_write                                        : std_logic;                     -- mm_interconnect_2:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	signal mm_interconnect_2_onchip_flash_0_data_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_2:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	signal mm_interconnect_2_onchip_flash_0_data_burstcount                                   : std_logic_vector(3 downto 0);  -- mm_interconnect_2:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	signal mm_interconnect_2_nios2_0_debug_mem_slave_readdata                                 : std_logic_vector(31 downto 0); -- nios2_0:debug_mem_slave_readdata -> mm_interconnect_2:nios2_0_debug_mem_slave_readdata
	signal mm_interconnect_2_nios2_0_debug_mem_slave_waitrequest                              : std_logic;                     -- nios2_0:debug_mem_slave_waitrequest -> mm_interconnect_2:nios2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_2_nios2_0_debug_mem_slave_debugaccess                              : std_logic;                     -- mm_interconnect_2:nios2_0_debug_mem_slave_debugaccess -> nios2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_2_nios2_0_debug_mem_slave_address                                  : std_logic_vector(8 downto 0);  -- mm_interconnect_2:nios2_0_debug_mem_slave_address -> nios2_0:debug_mem_slave_address
	signal mm_interconnect_2_nios2_0_debug_mem_slave_read                                     : std_logic;                     -- mm_interconnect_2:nios2_0_debug_mem_slave_read -> nios2_0:debug_mem_slave_read
	signal mm_interconnect_2_nios2_0_debug_mem_slave_byteenable                               : std_logic_vector(3 downto 0);  -- mm_interconnect_2:nios2_0_debug_mem_slave_byteenable -> nios2_0:debug_mem_slave_byteenable
	signal mm_interconnect_2_nios2_0_debug_mem_slave_write                                    : std_logic;                     -- mm_interconnect_2:nios2_0_debug_mem_slave_write -> nios2_0:debug_mem_slave_write
	signal mm_interconnect_2_nios2_0_debug_mem_slave_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_2:nios2_0_debug_mem_slave_writedata -> nios2_0:debug_mem_slave_writedata
	signal mm_interconnect_2_fifo_rx_in_csr_readdata                                          : std_logic_vector(31 downto 0); -- fifo_rx:wrclk_control_slave_readdata -> mm_interconnect_2:fifo_rx_in_csr_readdata
	signal mm_interconnect_2_fifo_rx_in_csr_address                                           : std_logic_vector(2 downto 0);  -- mm_interconnect_2:fifo_rx_in_csr_address -> fifo_rx:wrclk_control_slave_address
	signal mm_interconnect_2_fifo_rx_in_csr_read                                              : std_logic;                     -- mm_interconnect_2:fifo_rx_in_csr_read -> fifo_rx:wrclk_control_slave_read
	signal mm_interconnect_2_fifo_rx_in_csr_write                                             : std_logic;                     -- mm_interconnect_2:fifo_rx_in_csr_write -> fifo_rx:wrclk_control_slave_write
	signal mm_interconnect_2_fifo_rx_in_csr_writedata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_2:fifo_rx_in_csr_writedata -> fifo_rx:wrclk_control_slave_writedata
	signal mm_interconnect_2_altpll_0_pll_slave_readdata                                      : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_2:altpll_0_pll_slave_readdata
	signal mm_interconnect_2_altpll_0_pll_slave_address                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_2:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_2_altpll_0_pll_slave_read                                          : std_logic;                     -- mm_interconnect_2:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_2_altpll_0_pll_slave_write                                         : std_logic;                     -- mm_interconnect_2:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_2_altpll_0_pll_slave_writedata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_2:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_2_new_sdram_controller_0_s1_chipselect                             : std_logic;                     -- mm_interconnect_2:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	signal mm_interconnect_2_new_sdram_controller_0_s1_readdata                               : std_logic_vector(15 downto 0); -- new_sdram_controller_0:za_data -> mm_interconnect_2:new_sdram_controller_0_s1_readdata
	signal mm_interconnect_2_new_sdram_controller_0_s1_waitrequest                            : std_logic;                     -- new_sdram_controller_0:za_waitrequest -> mm_interconnect_2:new_sdram_controller_0_s1_waitrequest
	signal mm_interconnect_2_new_sdram_controller_0_s1_address                                : std_logic_vector(23 downto 0); -- mm_interconnect_2:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	signal mm_interconnect_2_new_sdram_controller_0_s1_read                                   : std_logic;                     -- mm_interconnect_2:new_sdram_controller_0_s1_read -> mm_interconnect_2_new_sdram_controller_0_s1_read:in
	signal mm_interconnect_2_new_sdram_controller_0_s1_byteenable                             : std_logic_vector(1 downto 0);  -- mm_interconnect_2:new_sdram_controller_0_s1_byteenable -> mm_interconnect_2_new_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_2_new_sdram_controller_0_s1_readdatavalid                          : std_logic;                     -- new_sdram_controller_0:za_valid -> mm_interconnect_2:new_sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_2_new_sdram_controller_0_s1_write                                  : std_logic;                     -- mm_interconnect_2:new_sdram_controller_0_s1_write -> mm_interconnect_2_new_sdram_controller_0_s1_write:in
	signal mm_interconnect_2_new_sdram_controller_0_s1_writedata                              : std_logic_vector(15 downto 0); -- mm_interconnect_2:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	signal mm_interconnect_2_sys_clk_timer_s1_chipselect                                      : std_logic;                     -- mm_interconnect_2:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_2_sys_clk_timer_s1_readdata                                        : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_2:sys_clk_timer_s1_readdata
	signal mm_interconnect_2_sys_clk_timer_s1_address                                         : std_logic_vector(2 downto 0);  -- mm_interconnect_2:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_2_sys_clk_timer_s1_write                                           : std_logic;                     -- mm_interconnect_2:sys_clk_timer_s1_write -> mm_interconnect_2_sys_clk_timer_s1_write:in
	signal mm_interconnect_2_sys_clk_timer_s1_writedata                                       : std_logic_vector(15 downto 0); -- mm_interconnect_2:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_2_pio_4_s1_chipselect                                              : std_logic;                     -- mm_interconnect_2:pio_4_s1_chipselect -> pio_4:chipselect
	signal mm_interconnect_2_pio_4_s1_readdata                                                : std_logic_vector(31 downto 0); -- pio_4:readdata -> mm_interconnect_2:pio_4_s1_readdata
	signal mm_interconnect_2_pio_4_s1_address                                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_2:pio_4_s1_address -> pio_4:address
	signal mm_interconnect_2_pio_4_s1_write                                                   : std_logic;                     -- mm_interconnect_2:pio_4_s1_write -> mm_interconnect_2_pio_4_s1_write:in
	signal mm_interconnect_2_pio_4_s1_writedata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_2:pio_4_s1_writedata -> pio_4:writedata
	signal mm_interconnect_2_pio_5_s1_chipselect                                              : std_logic;                     -- mm_interconnect_2:pio_5_s1_chipselect -> pio_5:chipselect
	signal mm_interconnect_2_pio_5_s1_readdata                                                : std_logic_vector(31 downto 0); -- pio_5:readdata -> mm_interconnect_2:pio_5_s1_readdata
	signal mm_interconnect_2_pio_5_s1_address                                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_2:pio_5_s1_address -> pio_5:address
	signal mm_interconnect_2_pio_5_s1_write                                                   : std_logic;                     -- mm_interconnect_2:pio_5_s1_write -> mm_interconnect_2_pio_5_s1_write:in
	signal mm_interconnect_2_pio_5_s1_writedata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_2:pio_5_s1_writedata -> pio_5:writedata
	signal mm_interconnect_2_pio_1_s1_chipselect                                              : std_logic;                     -- mm_interconnect_2:pio_1_s1_chipselect -> pio_1:chipselect
	signal mm_interconnect_2_pio_1_s1_readdata                                                : std_logic_vector(31 downto 0); -- pio_1:readdata -> mm_interconnect_2:pio_1_s1_readdata
	signal mm_interconnect_2_pio_1_s1_address                                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_2:pio_1_s1_address -> pio_1:address
	signal mm_interconnect_2_pio_1_s1_write                                                   : std_logic;                     -- mm_interconnect_2:pio_1_s1_write -> mm_interconnect_2_pio_1_s1_write:in
	signal mm_interconnect_2_pio_1_s1_writedata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_2:pio_1_s1_writedata -> pio_1:writedata
	signal mm_interconnect_2_pio_3_s1_readdata                                                : std_logic_vector(31 downto 0); -- pio_3:readdata -> mm_interconnect_2:pio_3_s1_readdata
	signal mm_interconnect_2_pio_3_s1_address                                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_2:pio_3_s1_address -> pio_3:address
	signal mm_interconnect_2_pio_6_s1_readdata                                                : std_logic_vector(31 downto 0); -- pio_6:readdata -> mm_interconnect_2:pio_6_s1_readdata
	signal mm_interconnect_2_pio_6_s1_address                                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_2:pio_6_s1_address -> pio_6:address
	signal mm_interconnect_2_uart_0_s1_chipselect                                             : std_logic;                     -- mm_interconnect_2:uart_0_s1_chipselect -> uart_0:chipselect
	signal mm_interconnect_2_uart_0_s1_readdata                                               : std_logic_vector(15 downto 0); -- uart_0:readdata -> mm_interconnect_2:uart_0_s1_readdata
	signal mm_interconnect_2_uart_0_s1_address                                                : std_logic_vector(2 downto 0);  -- mm_interconnect_2:uart_0_s1_address -> uart_0:address
	signal mm_interconnect_2_uart_0_s1_read                                                   : std_logic;                     -- mm_interconnect_2:uart_0_s1_read -> mm_interconnect_2_uart_0_s1_read:in
	signal mm_interconnect_2_uart_0_s1_begintransfer                                          : std_logic;                     -- mm_interconnect_2:uart_0_s1_begintransfer -> uart_0:begintransfer
	signal mm_interconnect_2_uart_0_s1_write                                                  : std_logic;                     -- mm_interconnect_2:uart_0_s1_write -> mm_interconnect_2_uart_0_s1_write:in
	signal mm_interconnect_2_uart_0_s1_writedata                                              : std_logic_vector(15 downto 0); -- mm_interconnect_2:uart_0_s1_writedata -> uart_0:writedata
	signal mm_interconnect_2_avalon_pwm_0_s1_readdata                                         : std_logic_vector(31 downto 0); -- avalon_pwm_0:avs_s1_readdata -> mm_interconnect_2:avalon_pwm_0_s1_readdata
	signal mm_interconnect_2_avalon_pwm_0_s1_address                                          : std_logic_vector(2 downto 0);  -- mm_interconnect_2:avalon_pwm_0_s1_address -> avalon_pwm_0:avs_s1_address
	signal mm_interconnect_2_avalon_pwm_0_s1_read                                             : std_logic;                     -- mm_interconnect_2:avalon_pwm_0_s1_read -> avalon_pwm_0:avs_s1_read
	signal mm_interconnect_2_avalon_pwm_0_s1_write                                            : std_logic;                     -- mm_interconnect_2:avalon_pwm_0_s1_write -> avalon_pwm_0:avs_s1_write
	signal mm_interconnect_2_avalon_pwm_0_s1_writedata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_2:avalon_pwm_0_s1_writedata -> avalon_pwm_0:avs_s1_writedata
	signal mm_interconnect_2_avalon_wb_s1_chipselect                                          : std_logic;                     -- mm_interconnect_2:avalon_wb_s1_chipselect -> avalon_wb:avs_s1_chipselect
	signal mm_interconnect_2_avalon_wb_s1_readdata                                            : std_logic_vector(31 downto 0); -- avalon_wb:avs_s1_readdata -> mm_interconnect_2:avalon_wb_s1_readdata
	signal mm_interconnect_2_avalon_wb_s1_waitrequest                                         : std_logic;                     -- avalon_wb:avs_s1_waitrequest -> mm_interconnect_2:avalon_wb_s1_waitrequest
	signal mm_interconnect_2_avalon_wb_s1_address                                             : std_logic_vector(7 downto 0);  -- mm_interconnect_2:avalon_wb_s1_address -> avalon_wb:avs_s1_address
	signal mm_interconnect_2_avalon_wb_s1_read                                                : std_logic;                     -- mm_interconnect_2:avalon_wb_s1_read -> avalon_wb:avs_s1_read
	signal mm_interconnect_2_avalon_wb_s1_byteenable                                          : std_logic_vector(3 downto 0);  -- mm_interconnect_2:avalon_wb_s1_byteenable -> avalon_wb:avs_s1_byteenable
	signal mm_interconnect_2_avalon_wb_s1_readdatavalid                                       : std_logic;                     -- avalon_wb:avs_s1_readdatavalid -> mm_interconnect_2:avalon_wb_s1_readdatavalid
	signal mm_interconnect_2_avalon_wb_s1_write                                               : std_logic;                     -- mm_interconnect_2:avalon_wb_s1_write -> avalon_wb:avs_s1_write
	signal mm_interconnect_2_avalon_wb_s1_writedata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_2:avalon_wb_s1_writedata -> avalon_wb:avs_s1_writedata
	signal mm_interconnect_2_timer_0_s1_chipselect                                            : std_logic;                     -- mm_interconnect_2:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_2_timer_0_s1_readdata                                              : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_2:timer_0_s1_readdata
	signal mm_interconnect_2_timer_0_s1_address                                               : std_logic_vector(2 downto 0);  -- mm_interconnect_2:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_2_timer_0_s1_write                                                 : std_logic;                     -- mm_interconnect_2:timer_0_s1_write -> mm_interconnect_2_timer_0_s1_write:in
	signal mm_interconnect_2_timer_0_s1_writedata                                             : std_logic_vector(15 downto 0); -- mm_interconnect_2:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_2_avalon_i2s_0_s1_address                                          : std_logic_vector(1 downto 0);  -- mm_interconnect_2:avalon_i2s_0_s1_address -> avalon_i2s_0:avs_s1_address
	signal mm_interconnect_2_avalon_i2s_0_s1_write                                            : std_logic;                     -- mm_interconnect_2:avalon_i2s_0_s1_write -> avalon_i2s_0:avs_s1_write
	signal mm_interconnect_2_avalon_i2s_0_s1_writedata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_2:avalon_i2s_0_s1_writedata -> avalon_i2s_0:avs_s1_writedata
	signal dma_rx_read_master_chipselect                                                      : std_logic;                     -- dma_rx:read_chipselect -> mm_interconnect_3:dma_rx_read_master_chipselect
	signal dma_rx_read_master_readdata                                                        : std_logic_vector(31 downto 0); -- mm_interconnect_3:dma_rx_read_master_readdata -> dma_rx:read_readdata
	signal dma_rx_read_master_waitrequest                                                     : std_logic;                     -- mm_interconnect_3:dma_rx_read_master_waitrequest -> dma_rx:read_waitrequest
	signal dma_rx_read_master_address                                                         : std_logic_vector(4 downto 0);  -- dma_rx:read_address -> mm_interconnect_3:dma_rx_read_master_address
	signal dma_rx_read_master_read                                                            : std_logic;                     -- dma_rx:read_read_n -> dma_rx_read_master_read:in
	signal dma_rx_read_master_readdatavalid                                                   : std_logic;                     -- mm_interconnect_3:dma_rx_read_master_readdatavalid -> dma_rx:read_readdatavalid
	signal mm_interconnect_3_fifo_rx_out_readdata                                             : std_logic_vector(31 downto 0); -- fifo_rx:avalonmm_read_slave_readdata -> mm_interconnect_3:fifo_rx_out_readdata
	signal mm_interconnect_3_fifo_rx_out_read                                                 : std_logic;                     -- mm_interconnect_3:fifo_rx_out_read -> fifo_rx:avalonmm_read_slave_read
	signal dma_tx_write_master_chipselect                                                     : std_logic;                     -- dma_tx:write_chipselect -> mm_interconnect_4:dma_tx_write_master_chipselect
	signal dma_tx_write_master_waitrequest                                                    : std_logic;                     -- mm_interconnect_4:dma_tx_write_master_waitrequest -> dma_tx:write_waitrequest
	signal dma_tx_write_master_address                                                        : std_logic_vector(4 downto 0);  -- dma_tx:write_address -> mm_interconnect_4:dma_tx_write_master_address
	signal dma_tx_write_master_byteenable                                                     : std_logic_vector(3 downto 0);  -- dma_tx:write_byteenable -> mm_interconnect_4:dma_tx_write_master_byteenable
	signal dma_tx_write_master_write                                                          : std_logic;                     -- dma_tx:write_write_n -> dma_tx_write_master_write:in
	signal dma_tx_write_master_writedata                                                      : std_logic_vector(31 downto 0); -- dma_tx:write_writedata -> mm_interconnect_4:dma_tx_write_master_writedata
	signal mm_interconnect_4_fifo_tx_in_write                                                 : std_logic;                     -- mm_interconnect_4:fifo_tx_in_write -> fifo_tx:avalonmm_write_slave_write
	signal mm_interconnect_4_fifo_tx_in_writedata                                             : std_logic_vector(31 downto 0); -- mm_interconnect_4:fifo_tx_in_writedata -> fifo_tx:avalonmm_write_slave_writedata
	signal irq_mapper_receiver0_irq                                                           : std_logic;                     -- fifo_rx:wrclk_control_slave_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                           : std_logic;                     -- jtaguart_0:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                           : std_logic;                     -- sys_clk_timer:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                           : std_logic;                     -- uart_0:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                           : std_logic;                     -- timer_0:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                                           : std_logic;                     -- dma_rx:dma_ctl_irq -> irq_mapper:receiver5_irq
	signal irq_mapper_receiver6_irq                                                           : std_logic;                     -- dma_tx:dma_ctl_irq -> irq_mapper:receiver6_irq
	signal vic_0_irq_input_irq                                                                : std_logic_vector(6 downto 0);  -- irq_mapper:sender_irq -> vic_0:irq_input_irq
	signal rst_controller_reset_out_reset                                                     : std_logic;                     -- rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_2:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal nios2_0_debug_reset_request_reset                                                  : std_logic;                     -- nios2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	signal rst_controller_001_reset_out_reset                                                 : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:avalon_i2s_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:avalon_i2s_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:avalon_i2s_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                                                 : std_logic;                     -- rst_controller_002:reset_out -> [irq_mapper:reset, mm_interconnect_0:fifo_rx_reset_in_reset_bridge_in_reset_reset, mm_interconnect_1:fifo_tx_reset_in_reset_bridge_in_reset_reset, mm_interconnect_2:intel_generic_serial_flash_interface_top_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:nios2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_3:dma_rx_reset_reset_bridge_in_reset_reset, mm_interconnect_4:dma_tx_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in, rst_translator:in_reset, vic_0:reset_reset]
	signal rst_controller_002_reset_out_reset_req                                             : std_logic;                     -- rst_controller_002:reset_req -> [nios2_0:reset_req, rst_translator:reset_req_in]
	signal rst_controller_003_reset_out_reset                                                 : std_logic;                     -- rst_controller_003:reset_out -> intel_generic_serial_flash_interface_top_0:reset_reset
	signal reset_reset_n_ports_inv                                                            : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal dma_tx_read_master_read_ports_inv                                                  : std_logic;                     -- dma_tx_read_master_read:inv -> mm_interconnect_2:dma_tx_read_master_read
	signal dma_rx_write_master_write_ports_inv                                                : std_logic;                     -- dma_rx_write_master_write:inv -> mm_interconnect_2:dma_rx_write_master_write
	signal mm_interconnect_2_jtaguart_0_avalon_jtag_slave_read_ports_inv                      : std_logic;                     -- mm_interconnect_2_jtaguart_0_avalon_jtag_slave_read:inv -> jtaguart_0:av_read_n
	signal mm_interconnect_2_jtaguart_0_avalon_jtag_slave_write_ports_inv                     : std_logic;                     -- mm_interconnect_2_jtaguart_0_avalon_jtag_slave_write:inv -> jtaguart_0:av_write_n
	signal mm_interconnect_2_dma_rx_control_port_slave_write_ports_inv                        : std_logic;                     -- mm_interconnect_2_dma_rx_control_port_slave_write:inv -> dma_rx:dma_ctl_write_n
	signal mm_interconnect_2_dma_tx_control_port_slave_write_ports_inv                        : std_logic;                     -- mm_interconnect_2_dma_tx_control_port_slave_write:inv -> dma_tx:dma_ctl_write_n
	signal mm_interconnect_2_new_sdram_controller_0_s1_read_ports_inv                         : std_logic;                     -- mm_interconnect_2_new_sdram_controller_0_s1_read:inv -> new_sdram_controller_0:az_rd_n
	signal mm_interconnect_2_new_sdram_controller_0_s1_byteenable_ports_inv                   : std_logic_vector(1 downto 0);  -- mm_interconnect_2_new_sdram_controller_0_s1_byteenable:inv -> new_sdram_controller_0:az_be_n
	signal mm_interconnect_2_new_sdram_controller_0_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_2_new_sdram_controller_0_s1_write:inv -> new_sdram_controller_0:az_wr_n
	signal mm_interconnect_2_sys_clk_timer_s1_write_ports_inv                                 : std_logic;                     -- mm_interconnect_2_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal mm_interconnect_2_pio_4_s1_write_ports_inv                                         : std_logic;                     -- mm_interconnect_2_pio_4_s1_write:inv -> pio_4:write_n
	signal mm_interconnect_2_pio_5_s1_write_ports_inv                                         : std_logic;                     -- mm_interconnect_2_pio_5_s1_write:inv -> pio_5:write_n
	signal mm_interconnect_2_pio_1_s1_write_ports_inv                                         : std_logic;                     -- mm_interconnect_2_pio_1_s1_write:inv -> pio_1:write_n
	signal mm_interconnect_2_uart_0_s1_read_ports_inv                                         : std_logic;                     -- mm_interconnect_2_uart_0_s1_read:inv -> uart_0:read_n
	signal mm_interconnect_2_uart_0_s1_write_ports_inv                                        : std_logic;                     -- mm_interconnect_2_uart_0_s1_write:inv -> uart_0:write_n
	signal mm_interconnect_2_timer_0_s1_write_ports_inv                                       : std_logic;                     -- mm_interconnect_2_timer_0_s1_write:inv -> timer_0:write_n
	signal dma_rx_read_master_read_ports_inv                                                  : std_logic;                     -- dma_rx_read_master_read:inv -> mm_interconnect_3:dma_rx_read_master_read
	signal dma_tx_write_master_write_ports_inv                                                : std_logic;                     -- dma_tx_write_master_write:inv -> mm_interconnect_4:dma_tx_write_master_write
	signal rst_controller_001_reset_out_reset_ports_inv                                       : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> avalon_i2s_0:csi_reset_n
	signal rst_controller_002_reset_out_reset_ports_inv                                       : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [avalon_pwm_0:csi_reset_n, avalon_wb:csi_reset_n, dma_rx:system_reset_n, dma_tx:system_reset_n, fifo_rx:reset_n, fifo_tx:reset_n, jtaguart_0:rst_n, new_sdram_controller_0:reset_n, nios2_0:reset_n, onchip_flash_0:reset_n, pio_1:reset_n, pio_3:reset_n, pio_4:reset_n, pio_5:reset_n, pio_6:reset_n, sys_clk_timer:reset_n, sysid:reset_n, timer_0:reset_n, uart_0:reset_n]

begin

	altpll_0 : component candy_gw_qsys_altpll_0
		port map (
			clk                => clk_clk,                                        --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,                 -- inclk_interface_reset.reset
			read               => mm_interconnect_2_altpll_0_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_2_altpll_0_pll_slave_write,     --                      .write
			address            => mm_interconnect_2_altpll_0_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_2_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_2_altpll_0_pll_slave_writedata, --                      .writedata
			c0                 => open,                                           --                    c0.clk
			c1                 => altpll_0_c1_clk,                                --                    c1.clk
			c2                 => sdclk_clk_clk,                                  --                    c2.clk
			c3                 => codec_clk_clk,                                  --                    c3.clk
			locked             => altpll_locked_export,                           --        locked_conduit.export
			scandone           => open,                                           --           (terminated)
			scandataout        => open,                                           --           (terminated)
			c4                 => open,                                           --           (terminated)
			areset             => '0',                                            --           (terminated)
			phasedone          => open,                                           --           (terminated)
			phasecounterselect => "000",                                          --           (terminated)
			phaseupdown        => '0',                                            --           (terminated)
			phasestep          => '0',                                            --           (terminated)
			scanclk            => '0',                                            --           (terminated)
			scanclkena         => '0',                                            --           (terminated)
			scandata           => '0',                                            --           (terminated)
			configupdate       => '0'                                             --           (terminated)
		);

	avalon_i2s_0 : component AVALON_I2S
		generic map (
			DATA_WIDTH => 32
		)
		port map (
			csi_reset_n        => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			avs_s1_address     => mm_interconnect_2_avalon_i2s_0_s1_address,    --                  s1.address
			avs_s1_write       => mm_interconnect_2_avalon_i2s_0_s1_write,      --                    .write
			avs_s1_writedata   => mm_interconnect_2_avalon_i2s_0_s1_writedata,  --                    .writedata
			LRCLK_I_MST        => i2s_lrclk_i_mst,                              -- external_connection.lrclk_i_mst
			DATA_I_MST         => i2s_data_i_mst,                               --                    .data_i_mst
			DATA_O_MST         => i2s_data_o_mst,                               --                    .data_o_mst
			LRCLK_O_SLV        => i2s_lrclk_o_slv,                              --                    .lrclk_o_slv
			DATA_O_SLV         => i2s_data_o_slv,                               --                    .data_o_slv
			BITCLK_O_SLV       => i2s_bitclk_o_slv,                             --                    .bitclk_o_slv
			av_mm2_address     => avalon_i2s_0_av_mm2_address,                  --              av_mm2.address
			av_mm2_waitrequest => avalon_i2s_0_av_mm2_waitrequest,              --                    .waitrequest
			av_mm2_read        => avalon_i2s_0_av_mm2_read,                     --                    .read
			av_mm2_readdata    => avalon_i2s_0_av_mm2_readdata,                 --                    .readdata
			av_mm1_address     => avalon_i2s_0_av_mm1_address,                  --              av_mm1.address
			av_mm1_write       => avalon_i2s_0_av_mm1_write,                    --                    .write
			av_mm1_writedata   => avalon_i2s_0_av_mm1_writedata,                --                    .writedata
			av_mm1_waitrequest => avalon_i2s_0_av_mm1_waitrequest,              --                    .waitrequest
			bit_clk_mst        => i2s_bclk_mst_clk                              --               clock.clk
		);

	avalon_pwm_0 : component AVALON2PWM
		generic map (
			WIDTH           => 3,
			PWM_COUNTER_MAX => 60000
		)
		port map (
			csi_clk          => altpll_0_c1_clk,                              --                 clk.clk
			csi_reset_n      => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			avs_s1_write     => mm_interconnect_2_avalon_pwm_0_s1_write,      --                  s1.write
			avs_s1_writedata => mm_interconnect_2_avalon_pwm_0_s1_writedata,  --                    .writedata
			avs_s1_address   => mm_interconnect_2_avalon_pwm_0_s1_address,    --                    .address
			avs_s1_read      => mm_interconnect_2_avalon_pwm_0_s1_read,       --                    .read
			avs_s1_readdata  => mm_interconnect_2_avalon_pwm_0_s1_readdata,   --                    .readdata
			PWM_OUT          => onbrd_led_pwm_out                             -- external_connection.pwm_out
		);

	avalon_wb : component AVALON2WB
		port map (
			avs_s1_address       => mm_interconnect_2_avalon_wb_s1_address,       --                  s1.address
			avs_s1_chipselect    => mm_interconnect_2_avalon_wb_s1_chipselect,    --                    .chipselect
			avs_s1_byteenable    => mm_interconnect_2_avalon_wb_s1_byteenable,    --                    .byteenable
			avs_s1_read          => mm_interconnect_2_avalon_wb_s1_read,          --                    .read
			avs_s1_write         => mm_interconnect_2_avalon_wb_s1_write,         --                    .write
			avs_s1_writedata     => mm_interconnect_2_avalon_wb_s1_writedata,     --                    .writedata
			avs_s1_waitrequest   => mm_interconnect_2_avalon_wb_s1_waitrequest,   --                    .waitrequest
			avs_s1_readdata      => mm_interconnect_2_avalon_wb_s1_readdata,      --                    .readdata
			avs_s1_readdatavalid => mm_interconnect_2_avalon_wb_s1_readdatavalid, --                    .readdatavalid
			ACK_I                => wb_ack_i,                                     -- external_connection.ack_i
			ADR_O                => wb_adr_o,                                     --                    .adr_o
			CLK_O                => wb_clk_o,                                     --                    .clk_o
			CYC_O                => wb_cyc_o,                                     --                    .cyc_o
			DAT_I                => wb_dat_i,                                     --                    .dat_i
			DAT_O                => wb_dat_o,                                     --                    .dat_o
			ERR_I                => wb_err_i,                                     --                    .err_i
			RST_O                => wb_rst_o,                                     --                    .rst_o
			RTY_I                => wb_rty_i,                                     --                    .rty_i
			SEL_O                => wb_sel_o,                                     --                    .sel_o
			STB_O                => wb_stb_o,                                     --                    .stb_o
			WE_O                 => wb_we_o,                                      --                    .we_o
			csi_reset_n          => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			csi_clk              => altpll_0_c1_clk                               --                 clk.clk
		);

	dma_rx : component candy_gw_qsys_dma_rx
		port map (
			clk                => altpll_0_c1_clk,                                             --                clk.clk
			system_reset_n     => rst_controller_002_reset_out_reset_ports_inv,                --              reset.reset_n
			dma_ctl_address    => mm_interconnect_2_dma_rx_control_port_slave_address,         -- control_port_slave.address
			dma_ctl_chipselect => mm_interconnect_2_dma_rx_control_port_slave_chipselect,      --                   .chipselect
			dma_ctl_readdata   => mm_interconnect_2_dma_rx_control_port_slave_readdata,        --                   .readdata
			dma_ctl_write_n    => mm_interconnect_2_dma_rx_control_port_slave_write_ports_inv, --                   .write_n
			dma_ctl_writedata  => mm_interconnect_2_dma_rx_control_port_slave_writedata,       --                   .writedata
			dma_ctl_irq        => irq_mapper_receiver5_irq,                                    --                irq.irq
			read_address       => dma_rx_read_master_address,                                  --        read_master.address
			read_chipselect    => dma_rx_read_master_chipselect,                               --                   .chipselect
			read_read_n        => dma_rx_read_master_read,                                     --                   .read_n
			read_readdata      => dma_rx_read_master_readdata,                                 --                   .readdata
			read_readdatavalid => dma_rx_read_master_readdatavalid,                            --                   .readdatavalid
			read_waitrequest   => dma_rx_read_master_waitrequest,                              --                   .waitrequest
			write_address      => dma_rx_write_master_address,                                 --       write_master.address
			write_chipselect   => dma_rx_write_master_chipselect,                              --                   .chipselect
			write_waitrequest  => dma_rx_write_master_waitrequest,                             --                   .waitrequest
			write_write_n      => dma_rx_write_master_write,                                   --                   .write_n
			write_writedata    => dma_rx_write_master_writedata,                               --                   .writedata
			write_byteenable   => dma_rx_write_master_byteenable                               --                   .byteenable
		);

	dma_tx : component candy_gw_qsys_dma_tx
		port map (
			clk                => altpll_0_c1_clk,                                             --                clk.clk
			system_reset_n     => rst_controller_002_reset_out_reset_ports_inv,                --              reset.reset_n
			dma_ctl_address    => mm_interconnect_2_dma_tx_control_port_slave_address,         -- control_port_slave.address
			dma_ctl_chipselect => mm_interconnect_2_dma_tx_control_port_slave_chipselect,      --                   .chipselect
			dma_ctl_readdata   => mm_interconnect_2_dma_tx_control_port_slave_readdata,        --                   .readdata
			dma_ctl_write_n    => mm_interconnect_2_dma_tx_control_port_slave_write_ports_inv, --                   .write_n
			dma_ctl_writedata  => mm_interconnect_2_dma_tx_control_port_slave_writedata,       --                   .writedata
			dma_ctl_irq        => irq_mapper_receiver6_irq,                                    --                irq.irq
			read_address       => dma_tx_read_master_address,                                  --        read_master.address
			read_chipselect    => dma_tx_read_master_chipselect,                               --                   .chipselect
			read_read_n        => dma_tx_read_master_read,                                     --                   .read_n
			read_readdata      => dma_tx_read_master_readdata,                                 --                   .readdata
			read_readdatavalid => dma_tx_read_master_readdatavalid,                            --                   .readdatavalid
			read_waitrequest   => dma_tx_read_master_waitrequest,                              --                   .waitrequest
			write_address      => dma_tx_write_master_address,                                 --       write_master.address
			write_chipselect   => dma_tx_write_master_chipselect,                              --                   .chipselect
			write_waitrequest  => dma_tx_write_master_waitrequest,                             --                   .waitrequest
			write_write_n      => dma_tx_write_master_write,                                   --                   .write_n
			write_writedata    => dma_tx_write_master_writedata,                               --                   .writedata
			write_byteenable   => dma_tx_write_master_byteenable                               --                   .byteenable
		);

	fifo_rx : component candy_gw_qsys_fifo_rx
		port map (
			wrclock                        => altpll_0_c1_clk,                              --   clk_in.clk
			reset_n                        => rst_controller_002_reset_out_reset_ports_inv, -- reset_in.reset_n
			avalonmm_write_slave_writedata => mm_interconnect_0_fifo_rx_in_writedata,       --       in.writedata
			avalonmm_write_slave_write     => mm_interconnect_0_fifo_rx_in_write,           --         .write
			avalonmm_read_slave_readdata   => mm_interconnect_3_fifo_rx_out_readdata,       --      out.readdata
			avalonmm_read_slave_read       => mm_interconnect_3_fifo_rx_out_read,           --         .read
			wrclk_control_slave_address    => mm_interconnect_2_fifo_rx_in_csr_address,     --   in_csr.address
			wrclk_control_slave_read       => mm_interconnect_2_fifo_rx_in_csr_read,        --         .read
			wrclk_control_slave_writedata  => mm_interconnect_2_fifo_rx_in_csr_writedata,   --         .writedata
			wrclk_control_slave_write      => mm_interconnect_2_fifo_rx_in_csr_write,       --         .write
			wrclk_control_slave_readdata   => mm_interconnect_2_fifo_rx_in_csr_readdata,    --         .readdata
			wrclk_control_slave_irq        => irq_mapper_receiver0_irq                      --   in_irq.irq
		);

	fifo_tx : component candy_gw_qsys_fifo_tx
		port map (
			wrclock                        => altpll_0_c1_clk,                              --   clk_in.clk
			reset_n                        => rst_controller_002_reset_out_reset_ports_inv, -- reset_in.reset_n
			avalonmm_write_slave_writedata => mm_interconnect_4_fifo_tx_in_writedata,       --       in.writedata
			avalonmm_write_slave_write     => mm_interconnect_4_fifo_tx_in_write,           --         .write
			avalonmm_read_slave_readdata   => mm_interconnect_1_fifo_tx_out_readdata,       --      out.readdata
			avalonmm_read_slave_read       => mm_interconnect_1_fifo_tx_out_read            --         .read
		);

	intel_generic_serial_flash_interface_top_0 : component candy_gw_qsys_intel_generic_serial_flash_interface_top_0
		generic map (
			DEVICE_FAMILY => "MAX 10",
			CHIP_SELS     => 1
		)
		port map (
			avl_csr_address       => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_address,       --   avl_csr.address
			avl_csr_read          => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_read,          --          .read
			avl_csr_readdata      => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_readdata,      --          .readdata
			avl_csr_write         => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_write,         --          .write
			avl_csr_writedata     => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_writedata,     --          .writedata
			avl_csr_waitrequest   => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest,   --          .waitrequest
			avl_csr_readdatavalid => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid, --          .readdatavalid
			avl_mem_write         => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_write,         --   avl_mem.write
			avl_mem_burstcount    => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_burstcount,    --          .burstcount
			avl_mem_waitrequest   => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest,   --          .waitrequest
			avl_mem_read          => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_read,          --          .read
			avl_mem_address       => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_address,       --          .address
			avl_mem_writedata     => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_writedata,     --          .writedata
			avl_mem_readdata      => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_readdata,      --          .readdata
			avl_mem_readdatavalid => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid, --          .readdatavalid
			avl_mem_byteenable    => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_byteenable,    --          .byteenable
			clk_clk               => altpll_0_c1_clk,                                                                    --       clk.clk
			reset_reset           => rst_controller_003_reset_out_reset,                                                 --     reset.reset
			qspi_pins_dclk        => qspi_dclk,                                                                          -- qspi_pins.dclk
			qspi_pins_ncs         => qspi_ncs,                                                                           --          .ncs
			qspi_pins_data        => qspi_data                                                                           --          .data
		);

	jtaguart_0 : component candy_gw_qsys_jtaguart_0
		port map (
			clk            => altpll_0_c1_clk,                                                --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                   --             reset.reset_n
			av_chipselect  => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                        --               irq.irq
		);

	new_sdram_controller_0 : component candy_gw_qsys_new_sdram_controller_0
		port map (
			clk            => altpll_0_c1_clk,                                                  --   clk.clk
			reset_n        => rst_controller_002_reset_out_reset_ports_inv,                     -- reset.reset_n
			az_addr        => mm_interconnect_2_new_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_2_new_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_2_new_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_2_new_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_2_new_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_2_new_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_2_new_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_2_new_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_2_new_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => new_sdram_controller_0_wire_addr,                                 --  wire.export
			zs_ba          => new_sdram_controller_0_wire_ba,                                   --      .export
			zs_cas_n       => new_sdram_controller_0_wire_cas_n,                                --      .export
			zs_cke         => new_sdram_controller_0_wire_cke,                                  --      .export
			zs_cs_n        => new_sdram_controller_0_wire_cs_n,                                 --      .export
			zs_dq          => new_sdram_controller_0_wire_dq,                                   --      .export
			zs_dqm         => new_sdram_controller_0_wire_dqm,                                  --      .export
			zs_ras_n       => new_sdram_controller_0_wire_ras_n,                                --      .export
			zs_we_n        => new_sdram_controller_0_wire_we_n                                  --      .export
		);

	nios2_0 : component candy_gw_qsys_nios2_0
		port map (
			clk                                 => altpll_0_c1_clk,                                       --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,                --                          .reset_req
			d_address                           => nios2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			eic_port_valid                      => vic_0_interrupt_controller_out_valid,                  --   interrupt_controller_in.valid
			eic_port_data                       => vic_0_interrupt_controller_out_data,                   --                          .data
			debug_reset_request                 => nios2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_2_nios2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_2_nios2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_2_nios2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_2_nios2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_2_nios2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_2_nios2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_2_nios2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_2_nios2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                   -- custom_instruction_master.readra
		);

	onchip_flash_0 : component altera_onchip_flash
		generic map (
			INIT_FILENAME                       => "",
			INIT_FILENAME_SIM                   => "",
			DEVICE_FAMILY                       => "MAX 10",
			PART_NAME                           => "10M16SAU169C8G",
			DEVICE_ID                           => "16",
			SECTOR1_START_ADDR                  => 0,
			SECTOR1_END_ADDR                    => 4095,
			SECTOR2_START_ADDR                  => 4096,
			SECTOR2_END_ADDR                    => 8191,
			SECTOR3_START_ADDR                  => 8192,
			SECTOR3_END_ADDR                    => 47103,
			SECTOR4_START_ADDR                  => 47104,
			SECTOR4_END_ADDR                    => 75775,
			SECTOR5_START_ADDR                  => 75776,
			SECTOR5_END_ADDR                    => 143359,
			MIN_VALID_ADDR                      => 0,
			MAX_VALID_ADDR                      => 143359,
			MIN_UFM_VALID_ADDR                  => 0,
			MAX_UFM_VALID_ADDR                  => 47103,
			SECTOR1_MAP                         => 1,
			SECTOR2_MAP                         => 2,
			SECTOR3_MAP                         => 3,
			SECTOR4_MAP                         => 4,
			SECTOR5_MAP                         => 5,
			ADDR_RANGE1_END_ADDR                => 143359,
			ADDR_RANGE2_END_ADDR                => 143359,
			ADDR_RANGE1_OFFSET                  => 1024,
			ADDR_RANGE2_OFFSET                  => 0,
			ADDR_RANGE3_OFFSET                  => 0,
			AVMM_DATA_ADDR_WIDTH                => 18,
			AVMM_DATA_DATA_WIDTH                => 32,
			AVMM_DATA_BURSTCOUNT_WIDTH          => 4,
			SECTOR_READ_PROTECTION_MODE         => 0,
			FLASH_SEQ_READ_DATA_COUNT           => 4,
			FLASH_ADDR_ALIGNMENT_BITS           => 2,
			FLASH_READ_CYCLE_MAX_INDEX          => 4,
			FLASH_RESET_CYCLE_MAX_INDEX         => 25,
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  => 120,
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX => 35000000,
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX => 30500,
			PARALLEL_MODE                       => true,
			READ_AND_WRITE_MODE                 => true,
			WRAPPING_BURST_MODE                 => false,
			IS_DUAL_BOOT                        => "False",
			IS_ERAM_SKIP                        => "True",
			IS_COMPRESSED_IMAGE                 => "False"
		)
		port map (
			clock                   => altpll_0_c1_clk,                                     --    clk.clk
			reset_n                 => rst_controller_002_reset_out_reset_ports_inv,        -- nreset.reset_n
			avmm_data_addr          => mm_interconnect_2_onchip_flash_0_data_address,       --   data.address
			avmm_data_read          => mm_interconnect_2_onchip_flash_0_data_read,          --       .read
			avmm_data_writedata     => mm_interconnect_2_onchip_flash_0_data_writedata,     --       .writedata
			avmm_data_write         => mm_interconnect_2_onchip_flash_0_data_write,         --       .write
			avmm_data_readdata      => mm_interconnect_2_onchip_flash_0_data_readdata,      --       .readdata
			avmm_data_waitrequest   => mm_interconnect_2_onchip_flash_0_data_waitrequest,   --       .waitrequest
			avmm_data_readdatavalid => mm_interconnect_2_onchip_flash_0_data_readdatavalid, --       .readdatavalid
			avmm_data_burstcount    => mm_interconnect_2_onchip_flash_0_data_burstcount,    --       .burstcount
			avmm_csr_addr           => mm_interconnect_2_onchip_flash_0_csr_address(0),     --    csr.address
			avmm_csr_read           => mm_interconnect_2_onchip_flash_0_csr_read,           --       .read
			avmm_csr_writedata      => mm_interconnect_2_onchip_flash_0_csr_writedata,      --       .writedata
			avmm_csr_write          => mm_interconnect_2_onchip_flash_0_csr_write,          --       .write
			avmm_csr_readdata       => mm_interconnect_2_onchip_flash_0_csr_readdata        --       .readdata
		);

	pio_1 : component candy_gw_qsys_pio_1
		port map (
			clk        => altpll_0_c1_clk,                              --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_2_pio_1_s1_address,           --                  s1.address
			write_n    => mm_interconnect_2_pio_1_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_2_pio_1_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_2_pio_1_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_2_pio_1_s1_readdata,          --                    .readdata
			in_port    => grove1_in_port,                               -- external_connection.export
			out_port   => grove1_out_port                               --                    .export
		);

	pio_3 : component candy_gw_qsys_pio_3
		port map (
			clk      => altpll_0_c1_clk,                              --                 clk.clk
			reset_n  => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_pio_3_s1_address,           --                  s1.address
			readdata => mm_interconnect_2_pio_3_s1_readdata,          --                    .readdata
			in_port  => pmod2_export                                  -- external_connection.export
		);

	pio_4 : component candy_gw_qsys_pio_4
		port map (
			clk        => altpll_0_c1_clk,                              --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_2_pio_4_s1_address,           --                  s1.address
			write_n    => mm_interconnect_2_pio_4_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_2_pio_4_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_2_pio_4_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_2_pio_4_s1_readdata,          --                    .readdata
			out_port   => codec_reset_export                            -- external_connection.export
		);

	pio_5 : component candy_gw_qsys_pio_4
		port map (
			clk        => altpll_0_c1_clk,                              --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_2_pio_5_s1_address,           --                  s1.address
			write_n    => mm_interconnect_2_pio_5_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_2_pio_5_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_2_pio_5_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_2_pio_5_s1_readdata,          --                    .readdata
			out_port   => oe_export                                     -- external_connection.export
		);

	pio_6 : component candy_gw_qsys_pio_6
		port map (
			clk      => altpll_0_c1_clk,                              --                 clk.clk
			reset_n  => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_pio_6_s1_address,           --                  s1.address
			readdata => mm_interconnect_2_pio_6_s1_readdata,          --                    .readdata
			in_port  => adc_export                                    -- external_connection.export
		);

	sys_clk_timer : component candy_gw_qsys_sys_clk_timer
		port map (
			clk        => altpll_0_c1_clk,                                    --   clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,       -- reset.reset_n
			address    => mm_interconnect_2_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_2_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_2_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_2_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_2_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                            --   irq.irq
		);

	sysid : component candy_gw_qsys_sysid
		port map (
			clock    => altpll_0_c1_clk,                                  --           clk.clk
			reset_n  => rst_controller_002_reset_out_reset_ports_inv,     --         reset.reset_n
			readdata => mm_interconnect_2_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_2_sysid_control_slave_address(0)  --              .address
		);

	timer_0 : component candy_gw_qsys_timer_0
		port map (
			clk        => altpll_0_c1_clk,                              --   clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_2_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_2_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_2_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_2_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_2_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver4_irq                      --   irq.irq
		);

	uart_0 : component candy_gw_qsys_uart_0
		port map (
			clk           => altpll_0_c1_clk,                              --                 clk.clk
			reset_n       => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address       => mm_interconnect_2_uart_0_s1_address,          --                  s1.address
			begintransfer => mm_interconnect_2_uart_0_s1_begintransfer,    --                    .begintransfer
			chipselect    => mm_interconnect_2_uart_0_s1_chipselect,       --                    .chipselect
			read_n        => mm_interconnect_2_uart_0_s1_read_ports_inv,   --                    .read_n
			write_n       => mm_interconnect_2_uart_0_s1_write_ports_inv,  --                    .write_n
			writedata     => mm_interconnect_2_uart_0_s1_writedata,        --                    .writedata
			readdata      => mm_interconnect_2_uart_0_s1_readdata,         --                    .readdata
			rxd           => uart_rxd,                                     -- external_connection.export
			txd           => uart_txd,                                     --                    .export
			cts_n         => uart_cts_n,                                   --                    .export
			rts_n         => uart_rts_n,                                   --                    .export
			irq           => irq_mapper_receiver3_irq                      --                 irq.irq
		);

	vic_0 : component candy_gw_qsys_vic_0
		port map (
			clk_clk                        => altpll_0_c1_clk,                              --                      clk.clk
			reset_reset                    => rst_controller_002_reset_out_reset,           --                    reset.reset
			irq_input_irq                  => vic_0_irq_input_irq,                          --                irq_input.irq
			csr_access_read                => mm_interconnect_2_vic_0_csr_access_read,      --               csr_access.read
			csr_access_write               => mm_interconnect_2_vic_0_csr_access_write,     --                         .write
			csr_access_address             => mm_interconnect_2_vic_0_csr_access_address,   --                         .address
			csr_access_writedata           => mm_interconnect_2_vic_0_csr_access_writedata, --                         .writedata
			csr_access_readdata            => mm_interconnect_2_vic_0_csr_access_readdata,  --                         .readdata
			interrupt_controller_out_valid => vic_0_interrupt_controller_out_valid,         -- interrupt_controller_out.valid
			interrupt_controller_out_data  => vic_0_interrupt_controller_out_data           --                         .data
		);

	mm_interconnect_0 : component candy_gw_qsys_mm_interconnect_0
		port map (
			altpll_0_c1_clk                                => altpll_0_c1_clk,                        --                              altpll_0_c1.clk
			clock_bridge_0_out_clk_clk                     => i2s_bclk_mst_clk,                       --                   clock_bridge_0_out_clk.clk
			avalon_i2s_0_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,     -- avalon_i2s_0_reset_reset_bridge_in_reset.reset
			fifo_rx_reset_in_reset_bridge_in_reset_reset   => rst_controller_002_reset_out_reset,     --   fifo_rx_reset_in_reset_bridge_in_reset.reset
			avalon_i2s_0_av_mm1_address                    => avalon_i2s_0_av_mm1_address,            --                      avalon_i2s_0_av_mm1.address
			avalon_i2s_0_av_mm1_waitrequest                => avalon_i2s_0_av_mm1_waitrequest,        --                                         .waitrequest
			avalon_i2s_0_av_mm1_write                      => avalon_i2s_0_av_mm1_write,              --                                         .write
			avalon_i2s_0_av_mm1_writedata                  => avalon_i2s_0_av_mm1_writedata,          --                                         .writedata
			fifo_rx_in_write                               => mm_interconnect_0_fifo_rx_in_write,     --                               fifo_rx_in.write
			fifo_rx_in_writedata                           => mm_interconnect_0_fifo_rx_in_writedata  --                                         .writedata
		);

	mm_interconnect_1 : component candy_gw_qsys_mm_interconnect_1
		port map (
			altpll_0_c1_clk                                => altpll_0_c1_clk,                        --                              altpll_0_c1.clk
			clock_bridge_0_out_clk_clk                     => i2s_bclk_mst_clk,                       --                   clock_bridge_0_out_clk.clk
			avalon_i2s_0_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,     -- avalon_i2s_0_reset_reset_bridge_in_reset.reset
			fifo_tx_reset_in_reset_bridge_in_reset_reset   => rst_controller_002_reset_out_reset,     --   fifo_tx_reset_in_reset_bridge_in_reset.reset
			avalon_i2s_0_av_mm2_address                    => avalon_i2s_0_av_mm2_address,            --                      avalon_i2s_0_av_mm2.address
			avalon_i2s_0_av_mm2_waitrequest                => avalon_i2s_0_av_mm2_waitrequest,        --                                         .waitrequest
			avalon_i2s_0_av_mm2_read                       => avalon_i2s_0_av_mm2_read,               --                                         .read
			avalon_i2s_0_av_mm2_readdata                   => avalon_i2s_0_av_mm2_readdata,           --                                         .readdata
			fifo_tx_out_read                               => mm_interconnect_1_fifo_tx_out_read,     --                              fifo_tx_out.read
			fifo_tx_out_readdata                           => mm_interconnect_1_fifo_tx_out_readdata  --                                         .readdata
		);

	mm_interconnect_2 : component candy_gw_qsys_mm_interconnect_2
		port map (
			altpll_0_c1_clk                                                              => altpll_0_c1_clk,                                                                    --                                                            altpll_0_c1.clk
			clk_0_clk_clk                                                                => clk_clk,                                                                            --                                                              clk_0_clk.clk
			clock_bridge_0_out_clk_clk                                                   => i2s_bclk_mst_clk,                                                                   --                                                 clock_bridge_0_out_clk.clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset                   => rst_controller_reset_out_reset,                                                     --                   altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			avalon_i2s_0_reset_reset_bridge_in_reset_reset                               => rst_controller_001_reset_out_reset,                                                 --                               avalon_i2s_0_reset_reset_bridge_in_reset.reset
			intel_generic_serial_flash_interface_top_0_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                                                 -- intel_generic_serial_flash_interface_top_0_reset_reset_bridge_in_reset.reset
			nios2_0_reset_reset_bridge_in_reset_reset                                    => rst_controller_002_reset_out_reset,                                                 --                                    nios2_0_reset_reset_bridge_in_reset.reset
			dma_rx_write_master_address                                                  => dma_rx_write_master_address,                                                        --                                                    dma_rx_write_master.address
			dma_rx_write_master_waitrequest                                              => dma_rx_write_master_waitrequest,                                                    --                                                                       .waitrequest
			dma_rx_write_master_byteenable                                               => dma_rx_write_master_byteenable,                                                     --                                                                       .byteenable
			dma_rx_write_master_chipselect                                               => dma_rx_write_master_chipselect,                                                     --                                                                       .chipselect
			dma_rx_write_master_write                                                    => dma_rx_write_master_write_ports_inv,                                                --                                                                       .write
			dma_rx_write_master_writedata                                                => dma_rx_write_master_writedata,                                                      --                                                                       .writedata
			dma_tx_read_master_address                                                   => dma_tx_read_master_address,                                                         --                                                     dma_tx_read_master.address
			dma_tx_read_master_waitrequest                                               => dma_tx_read_master_waitrequest,                                                     --                                                                       .waitrequest
			dma_tx_read_master_chipselect                                                => dma_tx_read_master_chipselect,                                                      --                                                                       .chipselect
			dma_tx_read_master_read                                                      => dma_tx_read_master_read_ports_inv,                                                  --                                                                       .read
			dma_tx_read_master_readdata                                                  => dma_tx_read_master_readdata,                                                        --                                                                       .readdata
			dma_tx_read_master_readdatavalid                                             => dma_tx_read_master_readdatavalid,                                                   --                                                                       .readdatavalid
			nios2_0_data_master_address                                                  => nios2_0_data_master_address,                                                        --                                                    nios2_0_data_master.address
			nios2_0_data_master_waitrequest                                              => nios2_0_data_master_waitrequest,                                                    --                                                                       .waitrequest
			nios2_0_data_master_byteenable                                               => nios2_0_data_master_byteenable,                                                     --                                                                       .byteenable
			nios2_0_data_master_read                                                     => nios2_0_data_master_read,                                                           --                                                                       .read
			nios2_0_data_master_readdata                                                 => nios2_0_data_master_readdata,                                                       --                                                                       .readdata
			nios2_0_data_master_readdatavalid                                            => nios2_0_data_master_readdatavalid,                                                  --                                                                       .readdatavalid
			nios2_0_data_master_write                                                    => nios2_0_data_master_write,                                                          --                                                                       .write
			nios2_0_data_master_writedata                                                => nios2_0_data_master_writedata,                                                      --                                                                       .writedata
			nios2_0_data_master_debugaccess                                              => nios2_0_data_master_debugaccess,                                                    --                                                                       .debugaccess
			nios2_0_instruction_master_address                                           => nios2_0_instruction_master_address,                                                 --                                             nios2_0_instruction_master.address
			nios2_0_instruction_master_waitrequest                                       => nios2_0_instruction_master_waitrequest,                                             --                                                                       .waitrequest
			nios2_0_instruction_master_read                                              => nios2_0_instruction_master_read,                                                    --                                                                       .read
			nios2_0_instruction_master_readdata                                          => nios2_0_instruction_master_readdata,                                                --                                                                       .readdata
			nios2_0_instruction_master_readdatavalid                                     => nios2_0_instruction_master_readdatavalid,                                           --                                                                       .readdatavalid
			altpll_0_pll_slave_address                                                   => mm_interconnect_2_altpll_0_pll_slave_address,                                       --                                                     altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                                     => mm_interconnect_2_altpll_0_pll_slave_write,                                         --                                                                       .write
			altpll_0_pll_slave_read                                                      => mm_interconnect_2_altpll_0_pll_slave_read,                                          --                                                                       .read
			altpll_0_pll_slave_readdata                                                  => mm_interconnect_2_altpll_0_pll_slave_readdata,                                      --                                                                       .readdata
			altpll_0_pll_slave_writedata                                                 => mm_interconnect_2_altpll_0_pll_slave_writedata,                                     --                                                                       .writedata
			avalon_i2s_0_s1_address                                                      => mm_interconnect_2_avalon_i2s_0_s1_address,                                          --                                                        avalon_i2s_0_s1.address
			avalon_i2s_0_s1_write                                                        => mm_interconnect_2_avalon_i2s_0_s1_write,                                            --                                                                       .write
			avalon_i2s_0_s1_writedata                                                    => mm_interconnect_2_avalon_i2s_0_s1_writedata,                                        --                                                                       .writedata
			avalon_pwm_0_s1_address                                                      => mm_interconnect_2_avalon_pwm_0_s1_address,                                          --                                                        avalon_pwm_0_s1.address
			avalon_pwm_0_s1_write                                                        => mm_interconnect_2_avalon_pwm_0_s1_write,                                            --                                                                       .write
			avalon_pwm_0_s1_read                                                         => mm_interconnect_2_avalon_pwm_0_s1_read,                                             --                                                                       .read
			avalon_pwm_0_s1_readdata                                                     => mm_interconnect_2_avalon_pwm_0_s1_readdata,                                         --                                                                       .readdata
			avalon_pwm_0_s1_writedata                                                    => mm_interconnect_2_avalon_pwm_0_s1_writedata,                                        --                                                                       .writedata
			avalon_wb_s1_address                                                         => mm_interconnect_2_avalon_wb_s1_address,                                             --                                                           avalon_wb_s1.address
			avalon_wb_s1_write                                                           => mm_interconnect_2_avalon_wb_s1_write,                                               --                                                                       .write
			avalon_wb_s1_read                                                            => mm_interconnect_2_avalon_wb_s1_read,                                                --                                                                       .read
			avalon_wb_s1_readdata                                                        => mm_interconnect_2_avalon_wb_s1_readdata,                                            --                                                                       .readdata
			avalon_wb_s1_writedata                                                       => mm_interconnect_2_avalon_wb_s1_writedata,                                           --                                                                       .writedata
			avalon_wb_s1_byteenable                                                      => mm_interconnect_2_avalon_wb_s1_byteenable,                                          --                                                                       .byteenable
			avalon_wb_s1_readdatavalid                                                   => mm_interconnect_2_avalon_wb_s1_readdatavalid,                                       --                                                                       .readdatavalid
			avalon_wb_s1_waitrequest                                                     => mm_interconnect_2_avalon_wb_s1_waitrequest,                                         --                                                                       .waitrequest
			avalon_wb_s1_chipselect                                                      => mm_interconnect_2_avalon_wb_s1_chipselect,                                          --                                                                       .chipselect
			dma_rx_control_port_slave_address                                            => mm_interconnect_2_dma_rx_control_port_slave_address,                                --                                              dma_rx_control_port_slave.address
			dma_rx_control_port_slave_write                                              => mm_interconnect_2_dma_rx_control_port_slave_write,                                  --                                                                       .write
			dma_rx_control_port_slave_readdata                                           => mm_interconnect_2_dma_rx_control_port_slave_readdata,                               --                                                                       .readdata
			dma_rx_control_port_slave_writedata                                          => mm_interconnect_2_dma_rx_control_port_slave_writedata,                              --                                                                       .writedata
			dma_rx_control_port_slave_chipselect                                         => mm_interconnect_2_dma_rx_control_port_slave_chipselect,                             --                                                                       .chipselect
			dma_tx_control_port_slave_address                                            => mm_interconnect_2_dma_tx_control_port_slave_address,                                --                                              dma_tx_control_port_slave.address
			dma_tx_control_port_slave_write                                              => mm_interconnect_2_dma_tx_control_port_slave_write,                                  --                                                                       .write
			dma_tx_control_port_slave_readdata                                           => mm_interconnect_2_dma_tx_control_port_slave_readdata,                               --                                                                       .readdata
			dma_tx_control_port_slave_writedata                                          => mm_interconnect_2_dma_tx_control_port_slave_writedata,                              --                                                                       .writedata
			dma_tx_control_port_slave_chipselect                                         => mm_interconnect_2_dma_tx_control_port_slave_chipselect,                             --                                                                       .chipselect
			fifo_rx_in_csr_address                                                       => mm_interconnect_2_fifo_rx_in_csr_address,                                           --                                                         fifo_rx_in_csr.address
			fifo_rx_in_csr_write                                                         => mm_interconnect_2_fifo_rx_in_csr_write,                                             --                                                                       .write
			fifo_rx_in_csr_read                                                          => mm_interconnect_2_fifo_rx_in_csr_read,                                              --                                                                       .read
			fifo_rx_in_csr_readdata                                                      => mm_interconnect_2_fifo_rx_in_csr_readdata,                                          --                                                                       .readdata
			fifo_rx_in_csr_writedata                                                     => mm_interconnect_2_fifo_rx_in_csr_writedata,                                         --                                                                       .writedata
			intel_generic_serial_flash_interface_top_0_avl_csr_address                   => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_address,       --                     intel_generic_serial_flash_interface_top_0_avl_csr.address
			intel_generic_serial_flash_interface_top_0_avl_csr_write                     => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_write,         --                                                                       .write
			intel_generic_serial_flash_interface_top_0_avl_csr_read                      => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_read,          --                                                                       .read
			intel_generic_serial_flash_interface_top_0_avl_csr_readdata                  => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_readdata,      --                                                                       .readdata
			intel_generic_serial_flash_interface_top_0_avl_csr_writedata                 => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_writedata,     --                                                                       .writedata
			intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid             => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid, --                                                                       .readdatavalid
			intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest               => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest,   --                                                                       .waitrequest
			intel_generic_serial_flash_interface_top_0_avl_mem_address                   => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_address,       --                     intel_generic_serial_flash_interface_top_0_avl_mem.address
			intel_generic_serial_flash_interface_top_0_avl_mem_write                     => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_write,         --                                                                       .write
			intel_generic_serial_flash_interface_top_0_avl_mem_read                      => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_read,          --                                                                       .read
			intel_generic_serial_flash_interface_top_0_avl_mem_readdata                  => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_readdata,      --                                                                       .readdata
			intel_generic_serial_flash_interface_top_0_avl_mem_writedata                 => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_writedata,     --                                                                       .writedata
			intel_generic_serial_flash_interface_top_0_avl_mem_burstcount                => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_burstcount,    --                                                                       .burstcount
			intel_generic_serial_flash_interface_top_0_avl_mem_byteenable                => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_byteenable,    --                                                                       .byteenable
			intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid             => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid, --                                                                       .readdatavalid
			intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest               => mm_interconnect_2_intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest,   --                                                                       .waitrequest
			jtaguart_0_avalon_jtag_slave_address                                         => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_address,                             --                                           jtaguart_0_avalon_jtag_slave.address
			jtaguart_0_avalon_jtag_slave_write                                           => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_write,                               --                                                                       .write
			jtaguart_0_avalon_jtag_slave_read                                            => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_read,                                --                                                                       .read
			jtaguart_0_avalon_jtag_slave_readdata                                        => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_readdata,                            --                                                                       .readdata
			jtaguart_0_avalon_jtag_slave_writedata                                       => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_writedata,                           --                                                                       .writedata
			jtaguart_0_avalon_jtag_slave_waitrequest                                     => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_waitrequest,                         --                                                                       .waitrequest
			jtaguart_0_avalon_jtag_slave_chipselect                                      => mm_interconnect_2_jtaguart_0_avalon_jtag_slave_chipselect,                          --                                                                       .chipselect
			new_sdram_controller_0_s1_address                                            => mm_interconnect_2_new_sdram_controller_0_s1_address,                                --                                              new_sdram_controller_0_s1.address
			new_sdram_controller_0_s1_write                                              => mm_interconnect_2_new_sdram_controller_0_s1_write,                                  --                                                                       .write
			new_sdram_controller_0_s1_read                                               => mm_interconnect_2_new_sdram_controller_0_s1_read,                                   --                                                                       .read
			new_sdram_controller_0_s1_readdata                                           => mm_interconnect_2_new_sdram_controller_0_s1_readdata,                               --                                                                       .readdata
			new_sdram_controller_0_s1_writedata                                          => mm_interconnect_2_new_sdram_controller_0_s1_writedata,                              --                                                                       .writedata
			new_sdram_controller_0_s1_byteenable                                         => mm_interconnect_2_new_sdram_controller_0_s1_byteenable,                             --                                                                       .byteenable
			new_sdram_controller_0_s1_readdatavalid                                      => mm_interconnect_2_new_sdram_controller_0_s1_readdatavalid,                          --                                                                       .readdatavalid
			new_sdram_controller_0_s1_waitrequest                                        => mm_interconnect_2_new_sdram_controller_0_s1_waitrequest,                            --                                                                       .waitrequest
			new_sdram_controller_0_s1_chipselect                                         => mm_interconnect_2_new_sdram_controller_0_s1_chipselect,                             --                                                                       .chipselect
			nios2_0_debug_mem_slave_address                                              => mm_interconnect_2_nios2_0_debug_mem_slave_address,                                  --                                                nios2_0_debug_mem_slave.address
			nios2_0_debug_mem_slave_write                                                => mm_interconnect_2_nios2_0_debug_mem_slave_write,                                    --                                                                       .write
			nios2_0_debug_mem_slave_read                                                 => mm_interconnect_2_nios2_0_debug_mem_slave_read,                                     --                                                                       .read
			nios2_0_debug_mem_slave_readdata                                             => mm_interconnect_2_nios2_0_debug_mem_slave_readdata,                                 --                                                                       .readdata
			nios2_0_debug_mem_slave_writedata                                            => mm_interconnect_2_nios2_0_debug_mem_slave_writedata,                                --                                                                       .writedata
			nios2_0_debug_mem_slave_byteenable                                           => mm_interconnect_2_nios2_0_debug_mem_slave_byteenable,                               --                                                                       .byteenable
			nios2_0_debug_mem_slave_waitrequest                                          => mm_interconnect_2_nios2_0_debug_mem_slave_waitrequest,                              --                                                                       .waitrequest
			nios2_0_debug_mem_slave_debugaccess                                          => mm_interconnect_2_nios2_0_debug_mem_slave_debugaccess,                              --                                                                       .debugaccess
			onchip_flash_0_csr_address                                                   => mm_interconnect_2_onchip_flash_0_csr_address,                                       --                                                     onchip_flash_0_csr.address
			onchip_flash_0_csr_write                                                     => mm_interconnect_2_onchip_flash_0_csr_write,                                         --                                                                       .write
			onchip_flash_0_csr_read                                                      => mm_interconnect_2_onchip_flash_0_csr_read,                                          --                                                                       .read
			onchip_flash_0_csr_readdata                                                  => mm_interconnect_2_onchip_flash_0_csr_readdata,                                      --                                                                       .readdata
			onchip_flash_0_csr_writedata                                                 => mm_interconnect_2_onchip_flash_0_csr_writedata,                                     --                                                                       .writedata
			onchip_flash_0_data_address                                                  => mm_interconnect_2_onchip_flash_0_data_address,                                      --                                                    onchip_flash_0_data.address
			onchip_flash_0_data_write                                                    => mm_interconnect_2_onchip_flash_0_data_write,                                        --                                                                       .write
			onchip_flash_0_data_read                                                     => mm_interconnect_2_onchip_flash_0_data_read,                                         --                                                                       .read
			onchip_flash_0_data_readdata                                                 => mm_interconnect_2_onchip_flash_0_data_readdata,                                     --                                                                       .readdata
			onchip_flash_0_data_writedata                                                => mm_interconnect_2_onchip_flash_0_data_writedata,                                    --                                                                       .writedata
			onchip_flash_0_data_burstcount                                               => mm_interconnect_2_onchip_flash_0_data_burstcount,                                   --                                                                       .burstcount
			onchip_flash_0_data_readdatavalid                                            => mm_interconnect_2_onchip_flash_0_data_readdatavalid,                                --                                                                       .readdatavalid
			onchip_flash_0_data_waitrequest                                              => mm_interconnect_2_onchip_flash_0_data_waitrequest,                                  --                                                                       .waitrequest
			pio_1_s1_address                                                             => mm_interconnect_2_pio_1_s1_address,                                                 --                                                               pio_1_s1.address
			pio_1_s1_write                                                               => mm_interconnect_2_pio_1_s1_write,                                                   --                                                                       .write
			pio_1_s1_readdata                                                            => mm_interconnect_2_pio_1_s1_readdata,                                                --                                                                       .readdata
			pio_1_s1_writedata                                                           => mm_interconnect_2_pio_1_s1_writedata,                                               --                                                                       .writedata
			pio_1_s1_chipselect                                                          => mm_interconnect_2_pio_1_s1_chipselect,                                              --                                                                       .chipselect
			pio_3_s1_address                                                             => mm_interconnect_2_pio_3_s1_address,                                                 --                                                               pio_3_s1.address
			pio_3_s1_readdata                                                            => mm_interconnect_2_pio_3_s1_readdata,                                                --                                                                       .readdata
			pio_4_s1_address                                                             => mm_interconnect_2_pio_4_s1_address,                                                 --                                                               pio_4_s1.address
			pio_4_s1_write                                                               => mm_interconnect_2_pio_4_s1_write,                                                   --                                                                       .write
			pio_4_s1_readdata                                                            => mm_interconnect_2_pio_4_s1_readdata,                                                --                                                                       .readdata
			pio_4_s1_writedata                                                           => mm_interconnect_2_pio_4_s1_writedata,                                               --                                                                       .writedata
			pio_4_s1_chipselect                                                          => mm_interconnect_2_pio_4_s1_chipselect,                                              --                                                                       .chipselect
			pio_5_s1_address                                                             => mm_interconnect_2_pio_5_s1_address,                                                 --                                                               pio_5_s1.address
			pio_5_s1_write                                                               => mm_interconnect_2_pio_5_s1_write,                                                   --                                                                       .write
			pio_5_s1_readdata                                                            => mm_interconnect_2_pio_5_s1_readdata,                                                --                                                                       .readdata
			pio_5_s1_writedata                                                           => mm_interconnect_2_pio_5_s1_writedata,                                               --                                                                       .writedata
			pio_5_s1_chipselect                                                          => mm_interconnect_2_pio_5_s1_chipselect,                                              --                                                                       .chipselect
			pio_6_s1_address                                                             => mm_interconnect_2_pio_6_s1_address,                                                 --                                                               pio_6_s1.address
			pio_6_s1_readdata                                                            => mm_interconnect_2_pio_6_s1_readdata,                                                --                                                                       .readdata
			sys_clk_timer_s1_address                                                     => mm_interconnect_2_sys_clk_timer_s1_address,                                         --                                                       sys_clk_timer_s1.address
			sys_clk_timer_s1_write                                                       => mm_interconnect_2_sys_clk_timer_s1_write,                                           --                                                                       .write
			sys_clk_timer_s1_readdata                                                    => mm_interconnect_2_sys_clk_timer_s1_readdata,                                        --                                                                       .readdata
			sys_clk_timer_s1_writedata                                                   => mm_interconnect_2_sys_clk_timer_s1_writedata,                                       --                                                                       .writedata
			sys_clk_timer_s1_chipselect                                                  => mm_interconnect_2_sys_clk_timer_s1_chipselect,                                      --                                                                       .chipselect
			sysid_control_slave_address                                                  => mm_interconnect_2_sysid_control_slave_address,                                      --                                                    sysid_control_slave.address
			sysid_control_slave_readdata                                                 => mm_interconnect_2_sysid_control_slave_readdata,                                     --                                                                       .readdata
			timer_0_s1_address                                                           => mm_interconnect_2_timer_0_s1_address,                                               --                                                             timer_0_s1.address
			timer_0_s1_write                                                             => mm_interconnect_2_timer_0_s1_write,                                                 --                                                                       .write
			timer_0_s1_readdata                                                          => mm_interconnect_2_timer_0_s1_readdata,                                              --                                                                       .readdata
			timer_0_s1_writedata                                                         => mm_interconnect_2_timer_0_s1_writedata,                                             --                                                                       .writedata
			timer_0_s1_chipselect                                                        => mm_interconnect_2_timer_0_s1_chipselect,                                            --                                                                       .chipselect
			uart_0_s1_address                                                            => mm_interconnect_2_uart_0_s1_address,                                                --                                                              uart_0_s1.address
			uart_0_s1_write                                                              => mm_interconnect_2_uart_0_s1_write,                                                  --                                                                       .write
			uart_0_s1_read                                                               => mm_interconnect_2_uart_0_s1_read,                                                   --                                                                       .read
			uart_0_s1_readdata                                                           => mm_interconnect_2_uart_0_s1_readdata,                                               --                                                                       .readdata
			uart_0_s1_writedata                                                          => mm_interconnect_2_uart_0_s1_writedata,                                              --                                                                       .writedata
			uart_0_s1_begintransfer                                                      => mm_interconnect_2_uart_0_s1_begintransfer,                                          --                                                                       .begintransfer
			uart_0_s1_chipselect                                                         => mm_interconnect_2_uart_0_s1_chipselect,                                             --                                                                       .chipselect
			vic_0_csr_access_address                                                     => mm_interconnect_2_vic_0_csr_access_address,                                         --                                                       vic_0_csr_access.address
			vic_0_csr_access_write                                                       => mm_interconnect_2_vic_0_csr_access_write,                                           --                                                                       .write
			vic_0_csr_access_read                                                        => mm_interconnect_2_vic_0_csr_access_read,                                            --                                                                       .read
			vic_0_csr_access_readdata                                                    => mm_interconnect_2_vic_0_csr_access_readdata,                                        --                                                                       .readdata
			vic_0_csr_access_writedata                                                   => mm_interconnect_2_vic_0_csr_access_writedata                                        --                                                                       .writedata
		);

	mm_interconnect_3 : component candy_gw_qsys_mm_interconnect_3
		port map (
			altpll_0_c1_clk                          => altpll_0_c1_clk,                        --                        altpll_0_c1.clk
			dma_rx_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,     -- dma_rx_reset_reset_bridge_in_reset.reset
			dma_rx_read_master_address               => dma_rx_read_master_address,             --                 dma_rx_read_master.address
			dma_rx_read_master_waitrequest           => dma_rx_read_master_waitrequest,         --                                   .waitrequest
			dma_rx_read_master_chipselect            => dma_rx_read_master_chipselect,          --                                   .chipselect
			dma_rx_read_master_read                  => dma_rx_read_master_read_ports_inv,      --                                   .read
			dma_rx_read_master_readdata              => dma_rx_read_master_readdata,            --                                   .readdata
			dma_rx_read_master_readdatavalid         => dma_rx_read_master_readdatavalid,       --                                   .readdatavalid
			fifo_rx_out_read                         => mm_interconnect_3_fifo_rx_out_read,     --                        fifo_rx_out.read
			fifo_rx_out_readdata                     => mm_interconnect_3_fifo_rx_out_readdata  --                                   .readdata
		);

	mm_interconnect_4 : component candy_gw_qsys_mm_interconnect_4
		port map (
			altpll_0_c1_clk                          => altpll_0_c1_clk,                        --                        altpll_0_c1.clk
			dma_tx_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,     -- dma_tx_reset_reset_bridge_in_reset.reset
			dma_tx_write_master_address              => dma_tx_write_master_address,            --                dma_tx_write_master.address
			dma_tx_write_master_waitrequest          => dma_tx_write_master_waitrequest,        --                                   .waitrequest
			dma_tx_write_master_byteenable           => dma_tx_write_master_byteenable,         --                                   .byteenable
			dma_tx_write_master_chipselect           => dma_tx_write_master_chipselect,         --                                   .chipselect
			dma_tx_write_master_write                => dma_tx_write_master_write_ports_inv,    --                                   .write
			dma_tx_write_master_writedata            => dma_tx_write_master_writedata,          --                                   .writedata
			fifo_tx_in_write                         => mm_interconnect_4_fifo_tx_in_write,     --                         fifo_tx_in.write
			fifo_tx_in_writedata                     => mm_interconnect_4_fifo_tx_in_writedata  --                                   .writedata
		);

	irq_mapper : component candy_gw_qsys_irq_mapper
		port map (
			clk           => altpll_0_c1_clk,                    --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			receiver6_irq => irq_mapper_receiver6_irq,           -- receiver6.irq
			sender_irq    => vic_0_irq_input_irq                 --    sender.irq
		);

	rst_controller : component candy_gw_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,           -- reset_in0.reset
			reset_in1      => nios2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                           --       clk.clk
			reset_out      => rst_controller_reset_out_reset,    -- reset_out.reset
			reset_req      => open,                              -- (terminated)
			reset_req_in0  => '0',                               -- (terminated)
			reset_req_in1  => '0',                               -- (terminated)
			reset_in2      => '0',                               -- (terminated)
			reset_req_in2  => '0',                               -- (terminated)
			reset_in3      => '0',                               -- (terminated)
			reset_req_in3  => '0',                               -- (terminated)
			reset_in4      => '0',                               -- (terminated)
			reset_req_in4  => '0',                               -- (terminated)
			reset_in5      => '0',                               -- (terminated)
			reset_req_in5  => '0',                               -- (terminated)
			reset_in6      => '0',                               -- (terminated)
			reset_req_in6  => '0',                               -- (terminated)
			reset_in7      => '0',                               -- (terminated)
			reset_req_in7  => '0',                               -- (terminated)
			reset_in8      => '0',                               -- (terminated)
			reset_req_in8  => '0',                               -- (terminated)
			reset_in9      => '0',                               -- (terminated)
			reset_req_in9  => '0',                               -- (terminated)
			reset_in10     => '0',                               -- (terminated)
			reset_req_in10 => '0',                               -- (terminated)
			reset_in11     => '0',                               -- (terminated)
			reset_req_in11 => '0',                               -- (terminated)
			reset_in12     => '0',                               -- (terminated)
			reset_req_in12 => '0',                               -- (terminated)
			reset_in13     => '0',                               -- (terminated)
			reset_req_in13 => '0',                               -- (terminated)
			reset_in14     => '0',                               -- (terminated)
			reset_req_in14 => '0',                               -- (terminated)
			reset_in15     => '0',                               -- (terminated)
			reset_req_in15 => '0'                                -- (terminated)
		);

	rst_controller_001 : component candy_gw_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios2_0_debug_reset_request_reset,  -- reset_in1.reset
			clk            => i2s_bclk_mst_clk,                   --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component candy_gw_qsys_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_0_debug_reset_request_reset,      -- reset_in1.reset
			clk            => altpll_0_c1_clk,                        --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_003 : component candy_gw_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios2_0_debug_reset_request_reset,  -- reset_in1.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	dma_tx_read_master_read_ports_inv <= not dma_tx_read_master_read;

	dma_rx_write_master_write_ports_inv <= not dma_rx_write_master_write;

	mm_interconnect_2_jtaguart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_2_jtaguart_0_avalon_jtag_slave_read;

	mm_interconnect_2_jtaguart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_2_jtaguart_0_avalon_jtag_slave_write;

	mm_interconnect_2_dma_rx_control_port_slave_write_ports_inv <= not mm_interconnect_2_dma_rx_control_port_slave_write;

	mm_interconnect_2_dma_tx_control_port_slave_write_ports_inv <= not mm_interconnect_2_dma_tx_control_port_slave_write;

	mm_interconnect_2_new_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_2_new_sdram_controller_0_s1_read;

	mm_interconnect_2_new_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_2_new_sdram_controller_0_s1_byteenable;

	mm_interconnect_2_new_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_2_new_sdram_controller_0_s1_write;

	mm_interconnect_2_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_2_sys_clk_timer_s1_write;

	mm_interconnect_2_pio_4_s1_write_ports_inv <= not mm_interconnect_2_pio_4_s1_write;

	mm_interconnect_2_pio_5_s1_write_ports_inv <= not mm_interconnect_2_pio_5_s1_write;

	mm_interconnect_2_pio_1_s1_write_ports_inv <= not mm_interconnect_2_pio_1_s1_write;

	mm_interconnect_2_uart_0_s1_read_ports_inv <= not mm_interconnect_2_uart_0_s1_read;

	mm_interconnect_2_uart_0_s1_write_ports_inv <= not mm_interconnect_2_uart_0_s1_write;

	mm_interconnect_2_timer_0_s1_write_ports_inv <= not mm_interconnect_2_timer_0_s1_write;

	dma_rx_read_master_read_ports_inv <= not dma_rx_read_master_read;

	dma_tx_write_master_write_ports_inv <= not dma_tx_write_master_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of candy_gw_qsys
